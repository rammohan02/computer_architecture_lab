// Half Adder module
module HA(in0, in1, sum, cout);
    input in0, in1;
    output sum, cout;

    assign sum=in0^in1;
    assign cout=in0&in1;

endmodule

// Full adder module
module FA (in0, in1, cin, sum, cout);
    input in0, in1, cin;
    output sum, cout;

    assign sum=in0^in1^cin;
    assign cout=(in0&in1)|((in0^in1)&cin);
endmodule

// module FA (input [105:0] x,input [105:0] y,input [105:0] z,output [105:0] u,output [105:0] v);
//     assign u = x^y^z;
//     assign v[0] = 0;
//     assign v[105:1] = (x&y) | (y&z) | (z&x);
// endmodule

// Module for multyplying mantessas
module MUL_MANT (ma, mb, pro);
    input[52:0]  ma, mb;
    output[52:0] pro;

    reg[52:0][52:0] pp;

    integer i;
    always @(*) begin
        for (i = 0; i<53; i++) begin
            pp[i] = ma&{53{mb[i]}};
            // if(mb[i]==1) begin
            //     pp[i] <= ma << i;
            // end
            // else begin
            //     pp[i] = 106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            // end
        end
    end

    // wire [105:0] u_l11, v_l11, u_l12, v_l12, u_l13, v_l13, u_l14, v_l14, u_l15, v_l15, u_l16, v_l16, u_l17, v_l17, u_l18, v_l18, u_l19, v_l19, u_l110, v_l110;

	// FA l11 (pp[0][105:0], pp[1][105:0], pp[2][105:0], u_l11[105:0], v_l11[105:0]);

    wire[2:1] s1, c1;
    wire[4:1] s2, c2;
    wire[6:1] s3, c3;
    wire[8:1] s4, c4;
    wire[10:1] s5, c5;
    wire[12:1] s6, c6;
    wire[14:1] s7, c7;
    wire[16:1] s8, c8;
    wire[18:1] s9, c9;
    wire[20:1] s10, c10;
    wire[22:1] s11, c11;
    wire[24:1] s12, c12;
    wire[26:1] s13, c13;
    wire[28:1] s14, c14;
    wire[30:1] s15, c15;
    wire[32:1] s16, c16;
    wire[34:1] s17, c17;
    wire[36:1] s18, c18;
    wire[38:1] s19, c19;
    wire[40:1] s20, c20;
    wire[42:1] s21, c21;
    wire[44:1] s22, c22;
    wire[46:1] s23, c23;
    wire[48:1] s24, c24;
    wire[50:1] s25, c25;
    wire[52:1] s26, c26;
    wire[54:1] s27, c27;
    wire[56:1] s28, c28;
    wire[58:1] s29, c29;
    wire[60:1] s30, c30;
    wire[62:1] s31, c31;
    wire[64:1] s32, c32;
    wire[66:1] s33, c33;
    wire[68:1] s34, c34;
    wire[70:1] s35, c35;
    wire[72:1] s36, c36;
    wire[74:1] s37, c37;
    wire[76:1] s38, c38;
    wire[78:1] s39, c39;
    wire[80:1] s40, c40;

    // 1
    HA ha1(pp[52][0], pp[51][1], s1[1], c1[1]);
    HA ha2(pp[51][2], pp[52][1], s1[2], c1[2]);

    // 2
    HA ha3(pp[50][1], pp[51][0], s2[1], c2[1]);
    FA fa1(pp[49][3], pp[50][2], s1[1], s2[2], c2[2]);
    FA fa2(pp[50][3], s1[2], c1[1], s2[3], c2[3]);
    FA fa4(pp[51][3], pp[52][2], c1[2], s2[4], c2[4]);

    // 3
    HA ha4(pp[49][1], pp[50][0], s3[1], c3[1]);
    FA fa5(pp[48][3], pp[49][2], s2[1], s3[2], c3[2]);
    FA fa6(pp[48][4], s2[2], c2[1], s3[3], c3[3]);
    FA fa7(pp[49][4], s2[3], c2[2], s3[4], c3[4]);
    FA fa8(pp[50][4], s2[4], c2[3], s3[5], c3[5]);
    FA fa9(pp[51][4], pp[52][3], c2[4], s3[6], c3[6]);

    // 4
    HA ha5(pp[48][1], pp[49][0], s4[1], c4[1]);
    FA fa10(pp[47][3], pp[48][2], s3[1], s4[2], c4[2]);
    FA fa11(pp[47][4], s3[2], c3[1], s4[3], c4[3]);
    FA fa12(pp[47][5], s3[3], c3[2], s4[4], c4[4]);
    FA fa13(pp[48][5], s3[4], c3[3], s4[5], c4[5]);
    FA fa14(pp[49][5], s3[5], c3[4], s4[6], c4[6]);
    FA fa15(pp[50][5], s3[6], c3[5], s4[7], c4[7]);
    FA fa16(pp[51][5], pp[52][4], c3[6], s4[8], c4[8]);

    // 5
    HA ha6(pp[47][1], pp[48][0], s5[1], c5[1]);
    FA fa17(pp[46][3], pp[47][2], s4[1], s5[2], c5[2]);
    FA fa18(pp[46][4], s4[2], c4[1], s5[3], c5[3]);
    FA fa19(pp[46][5], s4[3], c4[2], s5[4], c5[4]);
    FA fa20(pp[46][6], s4[4], c4[3], s5[5], c5[5]);
    FA fa21(pp[47][6], s4[5], c4[4], s5[6], c6[6]);
    FA fa22(pp[48][6], s4[6], c4[5], s5[7], c5[7]);
    FA fa23(pp[49][6], s4[7], c4[6], s5[8], c5[8]);
    FA fa24(pp[50][6], s4[8], c4[7], s5[9], c5[9]);
    FA fa25(pp[51][6], pp[52][5], c4[8], s5[10], c5[10]);

    // 6
    HA ha7(pp[46][1], pp[47][0], s6[1], c6[1]);
    FA fa26(pp[45][3], pp[46][2], s5[1], s6[2], c6[2]);
    FA fa27(pp[45][4], s5[2], c5[1], s6[3], c6[3]);
    FA fa28(pp[45][5], s5[3], c5[2], s6[4], c6[4]);
    FA fa29(pp[45][6], s5[4], c5[3], s6[5], c6[5]);
    FA fa30(pp[45][7], s5[5], c5[4], s6[6], c6[6]);
    FA fa31(pp[46][7], s5[6], c5[5], s6[7], c6[7]);
    FA fa32(pp[47][7], s5[7], c5[6], s6[8], c6[8]);
    FA fa33(pp[48][7], s5[8], c5[7], s6[9], c6[9]);
    FA fa34(pp[49][7], s5[9], c5[8], s6[10], c6[10]);
    FA fa35(pp[50][7], s5[10], c5[9], s6[11], c6[11]);
    FA fa36(pp[51][7], pp[52][6], c5[10], s6[12], c6[12]);

    // 7
    HA ha8(pp[45][1], pp[46][0], s7[1], c7[1]);
    FA fa37(pp[44][3], pp[45][2], s6[1], s7[2], c7[2]);
    FA fa38(pp[44][4], s6[2], c6[1], s7[3], c7[3]);
    FA fa39(pp[44][5], s6[3], c6[2], s7[4], c7[4]);
    FA fa40(pp[44][6], s6[4], c6[3], s7[5], c7[5]);
    FA fa41(pp[44][7], s6[5], c6[4], s7[6], c7[6]);
    FA fa42(pp[44][8], s6[6], c6[5], s7[7], c7[7]);
    FA fa43(pp[45][8], s6[7], c6[6], s7[8], c7[8]);
    FA fa44(pp[46][8], s6[8], c6[7], s7[9], c7[9]);
    FA fa45(pp[47][8], s6[9], c6[8], s7[10], c7[10]);
    FA fa46(pp[48][8], s6[10], c6[9], s7[11], c7[11]);
    FA fa47(pp[49][8], s6[11], c6[10], s7[12], c7[12]);
    FA fa48(pp[50][8], s6[12], c6[11], s7[13], c7[13]);
    FA fa49(pp[51][8], pp[52][7], c6[12], s7[14], c7[14]);

    // 8
    HA ha9(pp[44][1], pp[45][0], s8[1], c8[1]);
    FA fa50(pp[43][3], pp[44][2], s7[1], s8[2], c8[2]);
    FA fa51(pp[43][4], s7[2], c7[1], s8[3], c8[3]);
    FA fa52(pp[43][5], s7[3], c7[2], s8[4], c8[4]);
    FA fa53(pp[43][6], s7[4], c7[3], s8[5], c8[5]);
    FA fa54(pp[43][7], s7[5], c7[4], s8[6], c8[6]);
    FA fa55(pp[43][8], s7[6], c7[5], s8[7], c8[7]);
    FA fa56(pp[43][9], s7[7], c7[6], s8[8], c8[8]);
    FA fa57(pp[44][9], s7[8], c7[7], s8[9], c8[9]);
    FA fa58(pp[45][9], s7[9], c7[8], s8[10], c8[10]);
    FA fa59(pp[46][9], s7[10], c7[9], s8[11], c8[11]);
    FA fa60(pp[47][9], s7[11], c7[10], s8[12], c8[12]);
    FA fa61(pp[48][9], s7[12], c7[11], s8[13], c8[13]);
    FA fa62(pp[49][9], s7[13], c7[12], s8[14], c8[14]);
    FA fa63(pp[50][9], s7[14], c7[13], s8[15], c8[15]);
    FA fa64(pp[51][9], pp[52][8], c7[14], s8[16], c8[16]);

    // 9
    HA ha10(pp[43][1], pp[44][0], s9[1], c9[1]);
    FA fa65(pp[42][3], pp[43][2], s8[1], s9[2], c9[2]);
    FA fa66(pp[42][4], s8[2], c8[1], s9[3], c9[3]);
    FA fa67(pp[42][5], s8[3], c8[2], s9[4], c9[4]);
    FA fa68(pp[42][6], s8[4], c8[3], s9[5], c9[5]);
    FA fa69(pp[42][7], s8[5], c8[4], s9[6], c9[6]);
    FA fa70(pp[42][8], s8[6], c8[5], s9[7], c9[7]);
    FA fa71(pp[42][9], s8[7], c8[6], s9[8], c8[8]);
    FA fa72(pp[42][10], s8[8], c8[7], s9[9], c9[9]);
    FA fa73(pp[43][10], s8[9], c8[8], s9[10], c9[10]);
    FA fa74(pp[44][10], s8[10], c8[9], s9[11], c9[11]);
    FA fa75(pp[45][10], s8[11], c8[10], s9[12], c9[12]);
    FA fa76(pp[46][10], s8[12], c8[11], s9[13], c9[13]);
    FA fa77(pp[47][10], s8[13], c8[12], s9[14], c9[14]);
    FA fa78(pp[48][10], s8[14], c8[13], s9[15], c9[15]);
    FA fa79(pp[49][10], s8[15], c8[14], s9[16], c9[16]);
    FA fa80(pp[50][10], s8[16], c8[15], s9[17], c9[17]);
    FA fa81(pp[51][10], pp[52][9], c8[16], s9[18], c9[18]);

    // 10
    HA ha11(pp[41][1], pp[43][0], s10[1], c10[1]);
    FA fa82(pp[41][3], pp[42][2], s9[1], s10[2], c10[2]);
    FA fa83(pp[41][4], s9[2], c9[1], s10[3], c10[3]);
    FA fa84(pp[41][5], s9[3], c9[2], s10[4], c10[4]);
    FA fa85(pp[41][6], s9[4], c9[3], s10[5], c10[5]);
    FA fa86(pp[41][7], s9[5], c9[4], s10[6], c10[6]);
    FA fa87(pp[41][8], s9[6], c9[5], s10[7], c10[7]);
    FA fa88(pp[41][9], s9[7], c9[6], s10[8], c10[8]);
    FA fa89(pp[41][10], s9[8], c9[7], s10[9], c10[9]);
    FA fa90(pp[41][11], s9[9], c9[8], s10[10], c10[10]);
    FA fa91(pp[42][11], s9[10], c9[9], s10[11], c10[11]);
    FA fa92(pp[43][11], s9[11], c9[10], s10[12], c10[12]);
    FA fa93(pp[44][11], s9[12], c9[11], s10[13], c10[13]);
    FA fa94(pp[45][11], s9[13], c9[12], s10[14], c10[14]);
    FA fa95(pp[46][11], s9[14], c9[13], s10[15], c10[15]);
    FA fa96(pp[47][11], s9[15], c9[14], s10[16], c10[16]);
    FA fa97(pp[48][11], s9[16], c9[15], s10[17], c10[17]);
    FA fa98(pp[49][11], s9[17], c9[16], s10[18], c10[18]);
    FA fa99(pp[50][11], s9[18], c9[17], s10[19], c10[19]);
    FA fa100(pp[51][11], pp[52][10], c9[18], s10[20], c10[20]);

    // 11
    HA ha12(pp[41][1], pp[42][0], s11[1], c11[1]);
    FA fa101(pp[40][3], pp[41][2], s10[1], s11[2], c11[2]);
    FA fa102(pp[40][4], s10[2], c10[1], s11[3], c11[3]);
    FA fa103(pp[40][5], s10[3], c10[2], s11[4], c11[4]);
    FA fa104(pp[40][6], s10[4], c10[3], s11[5], c11[5]);
    FA fa105(pp[40][7], s10[5], c10[4], s11[6], c11[6]);
    FA fa106(pp[40][8], s10[6], c10[5], s11[7], c11[7]);
    FA fa107(pp[40][9], s10[7], c10[6], s11[8], c11[8]);
    FA fa108(pp[40][10], s10[8], c10[7], s11[9], c11[9]);
    FA fa109(pp[40][11], s10[9], c10[8], s11[10], c11[10]);
    FA fa110(pp[40][12], s10[10], c10[9], s11[11], c11[11]);
    FA fa111(pp[41][12], s10[11], c10[10], s11[12], c11[12]);
    FA fa112(pp[42][12], s10[12], c10[11], s11[13], c11[13]);
    FA fa113(pp[43][12], s10[13], c10[12], s11[14], c11[14]);
    FA fa114(pp[44][12], s10[14], c10[13], s11[15], c11[15]);
    FA fa115(pp[45][12], s10[15], c10[14], s11[16], c11[16]);
    FA fa116(pp[46][12], s10[16], c10[15], s11[17], c11[17]);
    FA fa117(pp[47][12], s10[17], c10[16], s11[18], c11[18]);
    FA fa118(pp[48][12], s10[18], c10[17], s11[19], c11[19]);
    FA fa119(pp[49][12], s10[19], c10[18], s11[20], c11[20]);
    FA fa120(pp[50][12], s10[20], c10[19], s11[21], c11[21]);
    FA fa121(pp[51][12], pp[52][11], c10[20], s11[22], c11[22]);

    // 12
    HA ha13(pp[40][1], pp[41][0], s12[1], c12[1]);
    FA fa122(pp[39][3], pp[40][2], s11[1], s12[2], c12[2]);
    FA fa123(pp[39][4], s11[2], c11[1], s12[3], c12[3]);
    FA fa124(pp[39][5], s11[3], c11[2], s12[4], c12[4]);
    FA fa125(pp[39][6], s11[4], c11[3], s12[5], c12[5]);
    FA fa126(pp[39][7], s11[5], c11[4], s12[6], c12[6]);
    FA fa127(pp[39][8], s11[6], c11[5], s12[7], c12[7]);
    FA fa128(pp[39][9], s11[7], c11[6], s12[8], c12[8]);
    FA fa129(pp[39][10], s11[8], c11[7], s12[9], c12[9]);
    FA fa130(pp[39][11], s11[9], c11[8], s12[10], c12[10]);
    FA fa131(pp[39][12], s11[10], c11[9], s12[11], c12[11]);
    FA fa132(pp[39][13], s11[11], c11[10], s12[12], c12[12]);
    FA fa133(pp[40][13], s11[12], c11[11], s12[13], c12[13]);
    FA fa134(pp[41][13], s11[13], c11[12], s12[14], c12[14]);
    FA fa135(pp[42][13], s11[14], c11[13], s12[15], c12[15]);
    FA fa136(pp[43][13], s11[15], c11[14], s12[16], c12[16]);
    FA fa137(pp[44][13], s11[16], c11[15], s12[17], c12[17]);
    FA fa138(pp[45][13], s11[17], c11[16], s12[18], c12[18]);
    FA fa139(pp[46][13], s11[18], c11[17], s12[19], c12[19]);
    FA fa140(pp[47][13], s11[19], c11[18], s12[20], c12[20]);
    FA fa141(pp[48][13], s11[20], c11[19], s12[21], c12[21]);
    FA fa142(pp[49][13], s11[21], c11[20], s12[22], c12[22]);
    FA fa143(pp[50][13], s11[22], c11[21], s12[23], c12[23]);
    FA fa144(pp[51][13], pp[52][12], c11[22], s12[24], c12[24]);

    // 13
    HA ha14(pp[39][1], pp[40][0], s13[1], c13[1]);
    FA fa145(pp[38][3], pp[39][2], s12[1], s13[2], c13[2]);
    FA fa146(pp[38][4], s12[2], c12[1], s13[3], c13[3]);
    FA fa147(pp[38][5], s12[3], c12[2], s13[4], c13[4]);
    FA fa148(pp[38][6], s12[4], c12[3], s13[5], c13[5]);
    FA fa149(pp[38][7], s12[5], c12[4], s13[6], c13[6]);
    FA fa150(pp[38][8], s12[6], c12[5], s13[7], c13[7]);
    FA fa151(pp[38][9], s12[7], c12[6], s13[8], c13[8]);
    FA fa152(pp[38][10], s12[8], c12[7], s13[9], c13[9]);
    FA fa153(pp[38][11], s12[9], c12[8], s13[10], c13[10]);
    FA fa154(pp[38][12], s12[10], c12[9], s13[11], c13[11]);
    FA fa155(pp[38][13], s12[11], c12[10], s13[12], c13[12]);
    FA fa156(pp[38][14], s12[12], c12[11], s13[13], c13[13]);
    FA fa157(pp[39][14], s12[13], c12[12], s13[14], c13[14]);
    FA fa158(pp[40][14], s12[14], c12[13], s13[15], c13[15]);
    FA fa159(pp[41][14], s12[15], c12[14], s13[16], c13[16]);
    FA fa160(pp[42][14], s12[16], c12[15], s13[17], c13[17]);
    FA fa161(pp[43][14], s12[17], c12[16], s13[18], c13[18]);
    FA fa162(pp[44][14], s12[18], c12[17], s13[19], c13[19]);
    FA fa163(pp[45][14], s12[19], c12[18], s13[20], c13[20]);
    FA fa164(pp[46][14], s12[20], c12[19], s13[21], c13[21]);
    FA fa165(pp[47][14], s12[21], c12[20], s13[22], c13[22]);
    FA fa166(pp[48][14], s12[22], c12[21], s13[23], c13[23]);
    FA fa167(pp[49][14], s12[23], c12[22], s13[24], c13[24]);
    FA fa168(pp[50][14], s12[24], c12[23], s13[25], c13[25]);
    FA fa169(pp[51][14], pp[52][13], c12[24], s13[26], c13[26]);

    // 14
    HA ha15(pp[38][1], pp[39][0], s14[1], c14[1]);
    FA fa170(pp[37][3], pp[38][2], s13[1], s14[2], c14[2]);
    FA fa171(pp[37][4], s13[2], c13[1], s14[3], c14[3]);
    FA fa172(pp[37][5], s13[3], c13[2], s14[4], c14[4]);
    FA fa173(pp[37][6], s13[4], c13[3], s14[5], c14[5]);
    FA fa174(pp[37][7], s13[5], c13[4], s14[6], c14[6]);
    FA fa175(pp[37][8], s13[6], c13[5], s14[7], c14[7]);
    FA fa176(pp[37][9], s13[7], c13[6], s14[8], c14[8]);
    FA fa177(pp[37][10], s13[8], c13[7], s14[9], c14[9]);
    FA fa178(pp[37][11], s13[9], c13[8], s14[10], c14[10]);
    FA fa179(pp[37][12], s13[10], c13[9], s14[11], c14[11]);
    FA fa180(pp[37][13], s13[11], c13[10], s14[12], c14[12]);
    FA fa181(pp[37][14], s13[12], c13[11], s14[13], c14[13]);
    FA fa182(pp[37][15], s13[13], c13[12], s14[14], c14[14]);
    FA fa183(pp[38][15], s13[14], c13[13], s14[15], c14[15]);
    FA fa184(pp[39][15], s13[15], c13[14], s14[16], c14[16]);
    FA fa185(pp[40][15], s13[16], c13[15], s14[17], c14[17]);
    FA fa186(pp[40][15], s13[17], c13[16], s14[18], c14[18]);
    FA fa187(pp[42][15], s13[18], c13[17], s14[19], c14[18]);
    FA fa188(pp[43][15], s13[19], c13[18], s14[20], c14[20]);
    FA fa189(pp[44][15], s13[20], c13[19], s14[21], c14[21]);
    FA fa190(pp[45][15], s13[21], c13[20], s14[22], c14[22]);
    FA fa191(pp[46][15], s13[22], c13[21], s14[23], c14[23]);
    FA fa192(pp[47][15], s13[23], c13[22], s14[24], c14[24]);
    FA fa193(pp[48][15], s13[24], c13[23], s14[25], c14[25]);
    FA fa194(pp[49][15], s13[25], c13[24], s14[26], c14[26]);
    FA fa195(pp[50][15], s13[26], c13[25], s14[27], c14[27]);
    FA fa196(pp[51][15], pp[52][14], c13[26], s14[28], c14[28]);


    // 15
    HA ha16(pp[37][1], pp[38][0], s15[1], c15[1]);
    FA fa197(pp[36][3], pp[37][2], s14[1], s15[2], c15[2]);
    FA fa198(pp[36][4], s14[2], c14[1], s15[3], c15[3]);
    FA fa199(pp[36][5], s14[3], c14[2], s15[4], c15[4]);
    FA fa200(pp[36][6], s14[4], c14[3], s15[5], c15[5]);
    FA fa201(pp[36][7], s14[5], c14[4], s15[6], c15[6]);
    FA fa202(pp[36][8], s14[6], c14[5], s15[7], c15[7]);
    FA fa203(pp[36][9], s14[7], c14[6], s15[8], c15[8]);
    FA fa204(pp[36][10], s14[8], c14[7], s15[9], c15[9]);
    FA fa205(pp[36][11], s14[9], c14[8], s15[10], c15[10]);
    FA fa206(pp[36][12], s14[10], c14[9], s15[11], c15[11]);
    FA fa207(pp[36][13], s14[11], c14[10], s15[12], c15[12]);
    FA fa208(pp[36][14], s14[12], c14[11], s15[13], c15[13]);
    FA fa209(pp[36][15], s14[13], c14[12], s15[14], c15[14]);
    FA fa210(pp[36][16], s14[14], c14[13], s15[15], c15[15]);
    FA fa211(pp[37][16], s14[15], c14[14], s15[16], c15[16]);
    FA fa212(pp[38][16], s14[16], c14[15], s15[17], c15[17]);
    FA fa213(pp[39][16], s14[17], c14[16], s15[18], c15[18]);
    FA fa214(pp[40][16], s14[18], c14[17], s15[19], c15[19]);
    FA fa215(pp[41][16], s14[19], c14[18], s15[20], c15[20]);
    FA fa216(pp[42][16], s14[20], c14[19], s15[21], c15[21]);
    FA fa217(pp[43][16], s14[21], c14[20], s15[22], c15[22]);
    FA fa218(pp[44][16], s14[22], c14[21], s15[23], c15[23]);
    FA fa219(pp[45][16], s14[23], c14[22], s15[24], c15[24]);
    FA fa220(pp[46][16], s14[24], c14[23], s15[25], c15[25]);
    FA fa221(pp[47][16], s14[25], c14[24], s15[26], c15[26]);
    FA fa222(pp[48][16], s14[26], c14[25], s15[27], c15[27]);
    FA fa223(pp[49][16], s14[27], c14[26], s15[28], c15[28]);
    FA fa224(pp[50][16], s14[28], c14[27], s15[29], c15[29]);
    FA fa225(pp[51][16], pp[52][15], c14[28], s15[30], c15[30]);

    // 16
    HA ha17(pp[36][1], pp[37][0], s16[1], c16[1]);
    FA fa226(pp[35][3], pp[36][2], s15[1], s16[2], c16[2]);
    FA fa227(pp[35][4], s15[2], c15[1], s16[3], c16[3]);
    FA fa228(pp[35][5], s15[3], c15[2], s16[4], c16[4]);
    FA fa229(pp[35][6], s15[4], c15[3], s16[5], c16[5]);
    FA fa230(pp[35][7], s15[5], c15[4], s16[6], c16[6]);
    FA fa231(pp[35][8], s15[6], c15[5], s16[7], c16[7]);
    FA fa232(pp[35][9], s15[7], c15[6], s16[8], c16[8]);
    FA fa233(pp[35][10], s15[8], c15[7], s16[9], c16[9]);
    FA fa234(pp[35][11], s15[9], c15[8], s16[10], c16[10]);
    FA fa235(pp[35][12], s15[10], c15[9], s16[11], c16[11]);
    FA fa236(pp[35][13], s15[11], c15[10], s16[12], c16[12]);
    FA fa237(pp[35][14], s15[12], c15[11], s16[13], c16[13]);
    FA fa238(pp[35][15], s15[13], c15[12], s16[14], c16[14]);
    FA fa239(pp[35][16], s15[14], c15[13], s16[15], c16[15]);
    FA fa240(pp[35][17], s15[15], c15[14], s16[16], c16[16]);
    FA fa241(pp[36][17], s15[16], c15[15], s16[17], c16[17]);
    FA fa242(pp[37][17], s15[17], c15[16], s16[18], c16[18]);
    FA fa243(pp[38][17], s15[18], c15[17], s16[19], c16[19]);
    FA fa244(pp[39][17], s15[19], c15[18], s16[20], c16[20]);
    FA fa245(pp[40][17], s15[20], c15[19], s16[21], c16[21]);
    FA fa246(pp[41][17], s15[21], c15[20], s16[22], c16[22]);
    FA fa247(pp[42][17], s15[22], c15[21], s16[23], c16[23]);
    FA fa248(pp[43][17], s15[23], c15[22], s16[24], c16[24]);
    FA fa249(pp[44][17], s15[24], c15[23], s16[25], c16[25]);
    FA fa250(pp[45][17], s15[25], c15[24], s16[26], c16[26]);
    FA fa251(pp[46][17], s15[26], c15[25], s16[27], c16[27]);
    FA fa252(pp[47][17], s15[27], c15[26], s16[28], c16[28]);
    FA fa253(pp[48][17], s15[28], c15[27], s16[29], c16[29]);
    FA fa254(pp[49][17], s15[29], c15[28], s16[30], c16[30]);
    FA fa255(pp[50][17], s15[30], c15[29], s16[31], c16[31]);
    FA fa256(pp[51][17], pp[52][16], c15[30], s16[32], c16[32]);

    // 17
    HA ha18(pp[35][1], pp[36][0], s17[1], c17[1]);
    FA fa257(pp[34][3], pp[35][2], s16[1], s17[2], c17[2]);
    FA fa258(pp[34][4], s16[2], c16[1], s17[3], c17[3]);
    FA fa259(pp[34][5], s16[3], c16[2], s17[4], c17[4]);
    FA fa260(pp[34][6], s16[4], c16[3], s17[5], c17[5]);
    FA fa261(pp[34][7], s16[5], c16[4], s17[6], c17[6]);
    FA fa262(pp[34][8], s16[6], c16[5], s17[7], c17[7]);
    FA fa263(pp[34][9], s16[7], c16[6], s17[8], c17[8]);
    FA fa264(pp[34][10], s16[8], c16[7], s17[9], c17[9]);
    FA fa265(pp[34][11], s16[9], c16[8], s17[10], c17[10]);
    FA fa266(pp[34][12], s16[10], c16[9], s17[11], c17[11]);
    FA fa267(pp[34][13], s16[11], c16[10], s17[12], c17[12]);
    FA fa268(pp[34][14], s16[12], c16[11], s17[13], c17[13]);
    FA fa269(pp[34][15], s16[13], c16[12], s17[14], c17[14]);
    FA fa270(pp[34][16], s16[14], c16[13], s17[15], c17[15]);
    FA fa271(pp[34][17], s16[15], c16[14], s17[16], c17[16]);
    FA fa272(pp[34][18], s16[16], c16[15], s17[17], c17[17]);
    FA fa273(pp[35][18], s16[17], c16[16], s17[18], c17[18]);
    FA fa274(pp[36][18], s16[18], c16[17], s17[19], c17[19]);
    FA fa275(pp[37][18], s16[19], c16[18], s17[20], c17[20]);
    FA fa276(pp[38][18], s16[20], c16[19], s17[21], c17[21]);
    FA fa277(pp[39][18], s16[21], c16[20], s17[22], c17[22]);
    FA fa278(pp[40][18], s16[22], c16[21], s17[23], c17[23]);
    FA fa279(pp[41][18], s16[23], c16[22], s17[24], c17[24]);
    FA fa280(pp[42][18], s16[24], c16[23], s17[25], c17[25]);
    FA fa281(pp[43][18], s16[25], c16[24], s17[26], c17[26]);
    FA fa282(pp[44][18], s16[26], c16[25], s17[27], c17[27]);
    FA fa283(pp[45][18], s16[27], c16[26], s17[28], c17[28]);
    FA fa284(pp[46][18], s16[28], c16[27], s17[29], c17[29]);
    FA fa285(pp[47][18], s16[29], c16[28], s17[30], c17[30]);
    FA fa286(pp[48][18], s16[30], c16[29], s17[31], c17[31]);
    FA fa287(pp[49][18], s16[31], c16[30], s17[32], c17[32]);
    FA fa288(pp[50][18], s16[31], c16[31], s17[33], c17[33]);
    FA fa289(pp[51][18], pp[52][17], c16[32], s17[34], c17[34]);

    // 18
    HA ha19(pp[34][1], pp[35][0], s18[1], c18[1]);
    FA fa290(pp[33][3], pp[34][2], s17[1], s18[2], c18[2]);
    FA fa291(pp[33][4], s17[2], c17[1], s18[3], c18[3]);
    FA fa292(pp[33][5], s17[3], c17[2], s18[4], c18[4]);
    FA fa293(pp[33][6], s17[4], c17[3], s18[5], c18[5]);
    FA fa294(pp[33][7], s17[5], c17[4], s18[6], c18[6]);
    FA fa295(pp[33][8], s17[6], c17[5], s18[7], c18[7]);
    FA fa296(pp[33][9], s17[7], c17[6], s18[8], c18[8]);
    FA fa297(pp[33][10], s17[8], c17[7], s18[9], c18[9]);
    FA fa298(pp[33][11], s17[9], c17[8], s18[10], c18[10]);
    FA fa299(pp[33][12], s17[10], c17[9], s18[11], c18[11]);
    FA fa300(pp[33][13], s17[11], c17[10], s18[12], c18[12]);
    FA fa301(pp[33][14], s17[12], c17[11], s18[13], c18[13]);
    FA fa302(pp[33][15], s17[13], c17[12], s18[14], c18[14]);
    FA fa303(pp[33][16], s17[14], c17[13], s18[15], c18[15]);
    FA fa304(pp[33][17], s17[15], c17[14], s18[16], c18[16]);
    FA fa305(pp[33][18], s17[16], c17[15], s18[17], c18[17]);
    FA fa306(pp[33][19], s17[17], c17[16], s18[18], c18[18]);
    FA fa307(pp[34][19], s17[18], c17[17], s18[19], c18[19]);
    FA fa308(pp[35][19], s17[19], c17[18], s18[20], c18[20]);
    FA fa309(pp[36][19], s17[20], c17[19], s18[21], c18[21]);
    FA fa310(pp[37][19], s17[21], c17[20], s18[22], c18[22]);
    FA fa311(pp[38][19], s17[22], c17[21], s18[23], c18[23]);
    FA fa312(pp[39][19], s17[23], c17[22], s18[24], c18[24]);
    FA fa313(pp[40][19], s17[24], c17[23], s18[25], c18[25]);
    FA fa314(pp[41][19], s17[25], c17[24], s18[26], c18[26]);
    FA fa315(pp[42][19], s17[26], c17[25], s18[27], c18[27]);
    FA fa316(pp[43][19], s17[27], c17[26], s18[28], c18[28]);
    FA fa317(pp[44][19], s17[28], c17[27], s18[29], c18[29]);
    FA fa318(pp[45][19], s17[29], c17[28], s18[30], c18[30]);
    FA fa319(pp[46][19], s17[30], c17[29], s18[31], c18[31]);
    FA fa320(pp[47][19], s17[31], c17[30], s18[32], c18[32]);
    FA fa321(pp[48][19], s17[32], c17[31], s18[33], c18[33]);
    FA fa322(pp[49][19], s17[33], c17[32], s18[34], c18[34]);
    FA fa323(pp[50][19], s17[34], c17[33], s18[35], c18[35]);
    FA fa324(pp[51][19], pp[52][18], c17[34], s18[36], c18[36]);

    // 19
    HA ha20(pp[33][1], pp[34][0], s19[1], c19[1]);
    FA fa325(pp[32][3], pp[33][2], s18[1], s19[2], c19[2]);
    FA fa326(pp[32][4], s18[2], c18[1], s19[3], c19[3]);
    FA fa327(pp[32][5], s18[3], c18[2], s19[4], c19[4]);
    FA fa328(pp[32][6], s18[4], c18[3], s19[5], c19[5]);
    FA fa329(pp[32][7], s18[5], c18[4], s19[6], c19[6]);
    FA fa330(pp[32][8], s18[6], c18[5], s19[7], c19[7]);
    FA fa331(pp[32][9], s18[7], c18[6], s19[8], c19[8]);
    FA fa332(pp[32][10], s18[8], c18[7], s19[9], c19[9]);
    FA fa333(pp[32][11], s18[9], c18[8], s19[10], c19[10]);
    FA fa334(pp[32][12], s18[10], c18[9], s19[11], c19[11]);
    FA fa335(pp[32][13], s18[11], c18[10], s19[12], c19[12]);
    FA fa336(pp[32][14], s18[12], c18[11], s19[13], c19[13]);
    FA fa337(pp[32][15], s18[13], c18[12], s19[14], c19[14]);
    FA fa338(pp[32][16], s18[14], c18[13], s19[15], c19[15]);
    FA fa339(pp[32][17], s18[15], c18[14], s19[16], c19[16]);
    FA fa340(pp[32][18], s18[16], c18[15], s19[17], c19[17]);
    FA fa341(pp[32][19], s18[17], c18[16], s19[18], c19[18]);
    FA fa342(pp[32][20], s18[18], c18[17], s19[19], c19[19]);
    FA fa343(pp[33][20], s18[19], c18[18], s19[20], c19[20]);
    FA fa344(pp[34][20], s18[20], c18[19], s19[21], c19[21]);
    FA fa345(pp[35][20], s18[21], c18[20], s19[22], c19[22]);
    FA fa346(pp[36][20], s18[22], c18[21], s19[23], c19[23]);
    FA fa347(pp[37][20], s18[23], c18[22], s19[24], c19[24]);
    FA fa348(pp[38][20], s18[24], c18[23], s19[25], c19[25]);
    FA fa349(pp[39][20], s18[25], c18[24], s19[26], c19[26]);
    FA fa350(pp[40][20], s18[26], c18[25], s19[27], c19[27]);
    FA fa351(pp[41][20], s18[27], c18[26], s19[28], c19[28]);
    FA fa352(pp[42][20], s18[28], c18[27], s19[29], c19[29]);
    FA fa353(pp[43][20], s18[29], c18[28], s19[30], c19[30]);
    FA fa354(pp[44][20], s18[30], c18[29], s19[31], c19[31]);
    FA fa355(pp[45][20], s18[31], c18[30], s19[32], c19[32]);
    FA fa356(pp[46][20], s18[32], c18[31], s19[33], c19[33]);
    FA fa357(pp[47][20], s18[33], c18[32], s19[34], c19[34]);
    FA fa358(pp[48][20], s18[34], c18[33], s19[35], c19[35]);
    FA fa359(pp[49][20], s18[35], c18[34], s19[36], c19[36]);
    FA fa360(pp[50][20], s18[36], c18[35], s19[37], c19[37]);
    FA fa361(pp[51][20], pp[52][19], c18[36], s19[38], c19[38]);

    // 20
    HA ha21(pp[32][1], pp[33][0], s20[1], c20[1]);
    FA fa362(pp[31][3], pp[32][2], s19[1], s20[2], c20[2]);
    FA fa363(pp[31][4], s19[2], c19[1], s20[3], c20[3]);
    FA fa364(pp[31][5], s19[3], c19[2], s20[4], c20[4]);
    FA fa365(pp[31][6], s19[4], c19[3], s20[5], c20[5]);
    FA fa366(pp[31][7], s19[5], c19[4], s20[6], c20[6]);
    FA fa367(pp[31][8], s19[6], c19[5], s20[7], c20[7]);
    FA fa368(pp[31][9], s19[7], c19[6], s20[8], c20[8]);
    FA fa369(pp[31][10], s19[8], c19[7], s20[9], c20[9]);
    FA fa370(pp[31][11], s19[9], c19[8], s20[10], c20[10]);
    FA fa371(pp[31][12], s19[10], c19[9], s20[11], c20[11]);
    FA fa372(pp[31][13], s19[11], c19[10], s20[12], c20[12]);
    FA fa373(pp[31][14], s19[12], c19[11], s20[13], c20[13]);
    FA fa374(pp[31][15], s19[13], c19[12], s20[14], c20[14]);
    FA fa375(pp[31][16], s19[14], c19[13], s20[15], c20[15]);
    FA fa376(pp[31][17], s19[15], c19[14], s20[16], c20[16]);
    FA fa377(pp[31][18], s19[16], c19[15], s20[17], c20[17]);
    FA fa378(pp[31][19], s19[17], c19[16], s20[18], c20[18]);
    FA fa379(pp[31][20], s19[18], c19[17], s20[19], c20[19]);
    FA fa380(pp[31][21], s19[19], c19[18], s20[20], c20[20]);
    FA fa381(pp[32][21], s19[20], c19[19], s20[21], c20[21]);
    FA fa382(pp[33][21], s19[21], c19[20], s20[22], c20[22]);
    FA fa383(pp[34][21], s19[22], c19[21], s20[23], c20[23]);
    FA fa384(pp[35][21], s19[23], c19[22], s20[24], c20[24]);
    FA fa385(pp[36][21], s19[24], c19[23], s20[25], c20[25]);
    FA fa386(pp[37][21], s19[25], c19[24], s20[26], c20[26]);
    FA fa387(pp[38][21], s19[26], c19[25], s20[27], c20[27]);
    FA fa388(pp[39][21], s19[27], c19[26], s20[28], c20[28]);
    FA fa389(pp[40][21], s19[28], c19[27], s20[29], c20[29]);
    FA fa390(pp[41][21], s19[29], c19[28], s20[30], c20[30]);
    FA fa391(pp[42][21], s19[30], c19[29], s20[31], c20[31]);
    FA fa392(pp[43][21], s19[31], c19[30], s20[32], c20[32]);
    FA fa393(pp[44][21], s19[32], c19[31], s20[33], c20[33]);
    FA fa394(pp[45][21], s19[33], c19[32], s20[34], c20[34]);
    FA fa395(pp[46][21], s19[34], c19[33], s20[35], c20[35]);
    FA fa396(pp[47][21], s19[35], c19[34], s20[36], c20[36]);
    FA fa397(pp[48][21], s19[36], c19[35], s20[37], c20[37]);
    FA fa398(pp[49][21], s19[37], c19[36], s20[38], c20[38]);
    FA fa399(pp[50][21], s19[38], c19[37], s20[39], c20[39]);
    FA fa400(pp[51][21], pp[52][20], c19[38], s20[40], c20[40]);

    // 21
    HA ha22(pp[31][1], pp[32][0], s21[1], c21[1]);
    FA fa401(pp[30][3], pp[31][2], s20[1], s21[2], c21[2]);
    FA fa402(pp[30][4], s20[2], c20[1], s21[3], s21[3]);
    FA fa403(pp[30][5], s20[3], c20[2], s21[4], s21[4]);
    FA fa404(pp[30][6], s20[4], c20[3], s21[5], s21[5]);
    FA fa405(pp[30][7], s20[5], c20[4], s21[6], s21[6]);
    FA fa406(pp[30][8], s20[6], c20[5], s21[7], s21[7]);
    FA fa407(pp[30][9], s20[7], c20[6], s21[8], s21[8]);
    FA fa408(pp[30][10], s20[8], c20[7], s21[9], s21[9]);
    FA fa409(pp[30][11], s20[9], c20[8], s21[10], s21[10]);
    FA fa410(pp[30][12], s20[10], c20[9], s21[11], s21[11]);
    FA fa411(pp[30][13], s20[11], c20[10], s21[12], s21[12]);
    FA fa412(pp[30][14], s20[12], c20[11], s21[13], s21[13]);
    FA fa413(pp[30][15], s20[13], c20[12], s21[14], s21[14]);
    FA fa414(pp[30][16], s20[14], c20[13], s21[15], s21[15]);
    FA fa415(pp[30][17], s20[15], c20[14], s21[16], s21[16]);
    FA fa416(pp[30][18], s20[16], c20[15], s21[17], s21[17]);
    FA fa417(pp[30][19], s20[17], c20[16], s21[18], s21[18]);
    FA fa418(pp[30][20], s20[18], c20[17], s21[19], s21[19]);
    FA fa419(pp[30][21], s20[19], c20[18], s21[20], s21[20]);
    FA fa420(pp[30][22], s20[20], c20[19], s21[21], s21[21]);
    FA fa421(pp[31][22], s20[21], c20[20], s21[22], s21[22]);
    FA fa422(pp[32][22], s20[22], c20[21], s21[23], s21[23]);
    FA fa423(pp[33][22], s20[23], c20[22], s21[23], s21[24]);
    FA fa424(pp[34][22], s20[24], c20[23], s21[25], s21[25]);
    FA fa425(pp[35][22], s20[25], c20[24], s21[26], s21[26]);
    FA fa426(pp[36][22], s20[26], c20[25], s21[27], s21[27]);
    FA fa427(pp[37][22], s20[27], c20[26], s21[28], s21[28]);
    FA fa428(pp[38][22], s20[28], c20[27], s21[29], s21[29]);
    FA fa429(pp[39][22], s20[29], c20[28], s21[30], s21[30]);
    FA fa430(pp[40][22], s20[30], c20[29], s21[31], s21[31]);
    FA fa431(pp[41][22], s20[31], c20[30], s21[32], s21[32]);
    FA fa432(pp[42][22], s20[32], c20[31], s21[33], s21[33]);
    FA fa433(pp[43][22], s20[33], c20[32], s21[34], s21[34]);
    FA fa434(pp[44][22], s20[34], c20[33], s21[35], s21[35]);
    FA fa435(pp[45][22], s20[35], c20[34], s21[36], s21[36]);
    FA fa436(pp[46][22], s20[36], c20[35], s21[37], s21[37]);
    FA fa437(pp[47][22], s20[37], c20[36], s21[38], s21[38]);
    FA fa438(pp[48][22], s20[38], c20[37], s21[39], s21[39]);
    FA fa439(pp[49][22], s20[39], c20[38], s21[40], s21[40]);
    FA fa440(pp[50][22], s20[40], c20[39], s21[41], s21[41]);
    FA fa441(pp[51][22], pp[52][21], c20[40], s21[42], s21[42]);

    // 22
    HA ha23(pp[30][1], pp[31][0], s22[2], c22[1]);
    FA fa442(pp[29][3], pp[30][2], s21[1], s22[2], c22[2]);
    FA fa443(pp[29][4], s21[2], c21[1], s22[3], c22[3]);
    FA fa444(pp[29][5], s21[3], c21[2], s22[4], c22[4]);
    FA fa445(pp[29][6], s21[4], c21[3], s22[5], c22[5]);
    FA fa446(pp[29][7], s21[5], c21[4], s22[6], c22[6]);
    FA fa447(pp[29][8], s21[6], c21[5], s22[7], c22[7]);
    FA fa448(pp[29][9], s21[7], c21[6], s22[8], c22[8]);
    FA fa449(pp[29][10], s21[8], c21[7], s22[9], c22[9]);
    FA fa450(pp[29][11], s21[9], c21[8], s22[10], c22[10]);
    FA fa451(pp[29][12], s21[10], c21[9], s22[11], c22[11]);
    FA fa452(pp[29][13], s21[11], c21[10], s22[12], c22[12]);
    FA fa453(pp[29][14], s21[12], c21[11], s22[13], c22[13]);
    FA fa454(pp[29][15], s21[13], c21[12], s22[14], c22[14]);
    FA fa455(pp[29][16], s21[14], c21[13], s22[15], c22[15]);
    FA fa456(pp[29][17], s21[15], c21[14], s22[16], c22[16]);
    FA fa457(pp[29][18], s21[16], c21[15], s22[17], c22[17]);
    FA fa458(pp[29][19], s21[17], c21[16], s22[18], c22[18]);
    FA fa459(pp[29][20], s21[18], c21[17], s22[19], c22[19]);
    FA fa460(pp[29][21], s21[19], c21[18], s22[20], c22[20]);
    FA fa461(pp[29][22], s21[20], c21[19], s22[21], c22[21]);
    FA fa462(pp[29][23], s21[21], c21[20], s22[22], c22[22]);
    FA fa463(pp[30][23], s21[22], c21[21], s22[23], c22[23]);
    FA fa464(pp[31][23], s21[23], c21[22], s22[24], c22[24]);
    FA fa465(pp[32][23], s21[24], c21[23], s22[25], c22[25]);
    FA fa466(pp[33][23], s21[25], c21[24], s22[26], c22[26]);
    FA fa467(pp[34][23], s21[26], c21[25], s22[27], c22[27]);
    FA fa468(pp[35][23], s21[27], c21[26], s22[28], c22[28]);
    FA fa469(pp[36][23], s21[28], c21[27], s22[29], c22[29]);
    FA fa470(pp[37][23], s21[29], c21[28], s22[30], c22[30]);
    FA fa471(pp[38][23], s21[30], c21[29], s22[31], c22[31]);
    FA fa472(pp[39][23], s21[31], c21[30], s22[32], c22[32]);
    FA fa473(pp[40][23], s21[32], c21[31], s22[33], c22[33]);
    FA fa474(pp[41][23], s21[33], c21[32], s22[34], c22[34]);
    FA fa475(pp[42][23], s21[34], c21[33], s22[35], c22[35]);
    FA fa476(pp[43][23], s21[35], c21[34], s22[36], c22[36]);
    FA fa477(pp[44][23], s21[36], c21[35], s22[37], c22[37]);
    FA fa478(pp[45][23], s21[37], c21[36], s22[38], c22[38]);
    FA fa479(pp[46][23], s21[38], c21[37], s22[39], c22[39]);
    FA fa480(pp[47][23], s21[39], c21[38], s22[40], c22[40]);
    FA fa481(pp[48][23], s21[40], c21[39], s22[41], c22[41]);
    FA fa482(pp[49][23], s21[41], c21[40], s22[42], c22[42]);
    FA fa483(pp[50][23], s21[42], c21[41], s22[43], c22[43]);
    FA fa484(pp[51][23], pp[52][22], c21[42], s22[44], c22[44]);

    // 23
    HA ha24(pp[29][1], pp[30][0], s23[1], c23[1]);
    FA fa485(pp[28][3], pp[29][2], s22[1], s23[2], c23[2]);
    FA fa486(pp[28][4], s22[2], c22[1], s23[3], c23[3]);
    FA fa487(pp[28][5], s22[3], c22[2], s23[4], c23[4]);
    FA fa488(pp[28][6], s22[4], c22[3], s23[5], c23[5]);
    FA fa489(pp[28][7], s22[5], c22[4], s23[6], c23[6]);
    FA fa490(pp[28][8], s22[6], c22[5], s23[7], c23[7]);
    FA fa491(pp[28][9], s22[7], c22[6], s23[8], c23[8]);
    FA fa492(pp[28][10], s22[8], c22[7], s23[9], c23[9]);
    FA fa493(pp[28][11], s22[9], c22[8], s23[10], c23[10]);
    FA fa494(pp[28][12], s22[10], c22[9], s23[11], c23[11]);
    FA fa495(pp[28][13], s22[11], c22[10], s23[12], c23[12]);
    FA fa496(pp[28][14], s22[12], c22[11], s23[13], c23[13]);
    FA fa497(pp[28][15], s22[13], c22[12], s23[14], c23[14]);
    FA fa498(pp[28][16], s22[14], c22[13], s23[15], c23[15]);
    FA fa499(pp[28][17], s22[15], c22[14], s23[16], c23[16]);
    FA fa500(pp[28][18], s22[16], c22[15], s23[17], c23[17]);
    FA fa501(pp[28][19], s22[17], c22[16], s23[18], c23[18]);
    FA fa502(pp[28][20], s22[18], c22[17], s23[19], c23[19]);
    FA fa503(pp[28][21], s22[19], c22[18], s23[20], c23[20]);
    FA fa504(pp[28][22], s22[20], c22[19], s23[21], c23[21]);
    FA fa505(pp[28][23], s22[21], c22[20], s23[22], c23[22]);
    FA fa506(pp[28][24], s22[22], c22[21], s23[23], c23[23]);
    FA fa507(pp[29][24], s22[23], c22[22], s23[24], c23[24]);
    FA fa508(pp[30][24], s22[24], c22[23], s23[25], c23[25]);
    FA fa509(pp[31][24], s22[25], c22[24], s23[26], c23[26]);
    FA fa510(pp[32][24], s22[26], c22[25], s23[27], c23[27]);
    FA fa511(pp[33][24], s22[27], c22[26], s23[28], c23[28]);
    FA fa512(pp[34][24], s22[28], c22[27], s23[29], c23[29]);
    FA fa513(pp[35][24], s22[29], c22[28], s23[30], c23[30]);
    FA fa514(pp[36][24], s22[30], c22[29], s23[31], c23[31]);
    FA fa515(pp[37][24], s22[31], c22[30], s23[32], c23[32]);
    FA fa516(pp[38][24], s22[32], c22[31], s23[33], c23[33]);
    FA fa517(pp[39][24], s22[33], c22[32], s23[34], c23[34]);
    FA fa518(pp[40][24], s22[34], c22[33], s23[35], c23[35]);
    FA fa519(pp[41][24], s22[35], c22[34], s23[36], c23[36]);
    FA fa520(pp[42][24], s22[36], c22[35], s23[37], c23[37]);
    FA fa521(pp[43][24], s22[37], c22[36], s23[38], c23[38]);
    FA fa522(pp[44][24], s22[38], c22[37], s23[39], c23[39]);
    FA fa523(pp[45][24], s22[39], c22[38], s23[40], c23[40]);
    FA fa524(pp[46][24], s22[40], c22[39], s23[41], c23[41]);
    FA fa525(pp[47][24], s22[41], c22[40], s23[42], c23[42]);
    FA fa526(pp[48][24], s22[42], c22[41], s23[43], c23[43]);
    FA fa527(pp[49][24], s22[43], c22[42], s23[44], c23[44]);
    FA fa528(pp[50][24], s22[44], c22[43], s23[45], c23[45]);
    FA fa529(pp[51][24], pp[52][23], c22[44], s23[46], c23[46]);

    // 24
    HA ha25(pp[28][1], pp[29][0], s24[1], c24[1]);
    FA fa530(pp[27][3], pp[28][2], s23[1], s24[2], c24[2]);
    FA fa531(pp[27][4], s23[2], c23[1], s24[3], c24[3]);
    FA fa532(pp[27][5], s23[3], c23[2], s24[4], c24[4]);
    FA fa533(pp[27][6], s23[4], c23[3], s24[5], c24[5]);
    FA fa534(pp[27][7], s23[5], c23[4], s24[6], c24[6]);
    FA fa535(pp[27][8], s23[6], c23[5], s24[7], c24[7]);
    FA fa536(pp[27][9], s23[7], c23[6], s24[8], c24[8]);
    FA fa537(pp[27][10], s23[8], c23[7], s24[9], c24[9]);
    FA fa538(pp[27][11], s23[9], c23[8], s24[10], c24[10]);
    FA fa539(pp[27][12], s23[10], c23[9], s24[11], c24[11]);
    FA fa540(pp[27][13], s23[11], c23[10], s24[12], c24[12]);
    FA fa541(pp[27][14], s23[12], c23[11], s24[13], c24[13]);
    FA fa542(pp[27][15], s23[13], c23[12], s24[14], c24[14]);
    FA fa543(pp[27][16], s23[14], c23[13], s24[15], c24[15]);
    FA fa544(pp[27][17], s23[15], c23[14], s24[16], c24[16]);
    FA fa545(pp[27][18], s23[16], c23[15], s24[17], c24[17]);
    FA fa546(pp[27][19], s23[17], c23[16], s24[18], c24[18]);
    FA fa547(pp[27][20], s23[18], c23[17], s24[19], c24[19]);
    FA fa548(pp[27][21], s23[19], c23[18], s24[20], c24[20]);
    FA fa549(pp[27][22], s23[20], c23[19], s24[21], c24[21]);
    FA fa550(pp[27][23], s23[21], c23[20], s24[22], c24[22]);
    FA fa551(pp[27][24], s23[22], c23[21], s24[23], c24[23]);
    FA fa552(pp[27][25], s23[23], c23[22], s24[24], c24[24]);
    FA fa553(pp[28][25], s23[24], c23[23], s24[25], c24[25]);
    FA fa554(pp[29][25], s23[25], c23[24], s24[26], c24[26]);
    FA fa555(pp[30][25], s23[26], c23[25], s24[27], c24[27]);
    FA fa556(pp[31][25], s23[27], c23[26], s24[28], c24[28]);
    FA fa557(pp[32][25], s23[28], c23[27], s24[29], c24[29]);
    FA fa558(pp[33][25], s23[29], c23[28], s24[30], c24[30]);
    FA fa559(pp[34][25], s23[30], c23[29], s24[31], c24[31]);
    FA fa560(pp[35][25], s23[31], c23[30], s24[32], c24[32]);
    FA fa561(pp[36][25], s23[32], c23[31], s24[33], c24[33]);
    FA fa562(pp[37][25], s23[33], c23[32], s24[34], c24[34]);
    FA fa563(pp[38][25], s23[34], c23[33], s24[35], c24[35]);
    FA fa564(pp[39][25], s23[35], c23[34], s24[36], c24[36]);
    FA fa565(pp[40][25], s23[36], c23[35], s24[37], c24[37]);
    FA fa566(pp[41][25], s23[37], c23[36], s24[38], c24[38]);
    FA fa567(pp[42][25], s23[38], c23[37], s24[39], c24[39]);
    FA fa568(pp[43][25], s23[39], c23[38], s24[40], c24[40]);
    FA fa569(pp[44][25], s23[40], c23[39], s24[41], c24[41]);
    FA fa570(pp[45][25], s23[41], c23[40], s24[42], c24[42]);
    FA fa571(pp[46][25], s23[42], c23[41], s24[43], c24[43]);
    FA fa572(pp[47][25], s23[43], c23[42], s24[44], c24[44]);
    FA fa573(pp[48][25], s23[44], c23[43], s24[45], c24[45]);
    FA fa574(pp[49][25], s23[45], c23[44], s24[46], c24[46]);
    FA fa575(pp[50][25], s23[46], c23[45], s24[47], c24[47]);
    FA fa576(pp[51][25], pp[52][24], c23[46], s24[48], c24[48]);

    // 25
    HA ha26(pp[27][1], pp[28][0], s25[1], c25[1]);
    FA fa577(pp[26][3], pp[27][2], s24[1], s25[2], c25[2]);
    FA fa578(pp[26][4], s24[2], c24[1], s25[3], c25[3]);
    FA fa579(pp[26][5], s24[3], c24[2], s25[4], c25[4]);
    FA fa580(pp[26][6], s24[4], c24[3], s25[5], c25[5]);
    FA fa581(pp[26][7], s24[5], c24[4], s25[6], c25[6]);
    FA fa582(pp[26][8], s24[6], c24[5], s25[7], c25[7]);
    FA fa583(pp[26][9], s24[7], c24[6], s25[8], c25[8]);
    FA fa584(pp[26][10], s24[8], c24[7], s25[9], c25[9]);
    FA fa585(pp[26][11], s24[9], c24[8], s25[10], c25[10]);
    FA fa586(pp[26][12], s24[10], c24[9], s25[11], c25[11]);
    FA fa587(pp[26][13], s24[11], c24[10], s25[12], c25[12]);
    FA fa588(pp[26][14], s24[12], c24[11], s25[13], c25[13]);
    FA fa589(pp[26][15], s24[13], c24[12], s25[14], c25[14]);
    FA fa590(pp[26][16], s24[14], c24[13], s25[15], c25[15]);
    FA fa591(pp[26][17], s24[15], c24[14], s25[16], c25[16]);
    FA fa592(pp[26][18], s24[16], c24[15], s25[17], c25[17]);
    FA fa593(pp[26][19], s24[17], c24[16], s25[18], c25[18]);
    FA fa594(pp[26][20], s24[18], c24[17], s25[19], c25[19]);
    FA fa595(pp[26][21], s24[19], c24[18], s25[20], c25[20]);
    FA fa596(pp[26][22], s24[20], c24[19], s25[21], c25[21]);
    FA fa597(pp[26][23], s24[21], c24[20], s25[22], c25[22]);
    FA fa598(pp[26][24], s24[22], c24[21], s25[23], c25[23]);
    FA fa599(pp[26][25], s24[23], c24[22], s25[24], c25[24]);
    FA fa600(pp[26][26], s24[24], c24[23], s25[25], c25[25]);
    FA fa601(pp[27][26], s24[25], c24[24], s25[26], c25[26]);
    FA fa602(pp[28][26], s24[26], c24[25], s25[27], c25[27]);
    FA fa603(pp[29][26], s24[27], c24[26], s25[28], c25[28]);
    FA fa604(pp[30][26], s24[28], c24[27], s25[29], c25[29]);
    FA fa605(pp[31][26], s24[29], c24[28], s25[30], c25[30]);
    FA fa606(pp[32][26], s24[30], c24[29], s25[31], c25[31]);
    FA fa607(pp[33][26], s24[31], c24[30], s25[32], c25[32]);
    FA fa608(pp[34][26], s24[32], c24[31], s25[33], c25[33]);
    FA fa609(pp[35][26], s24[33], c24[32], s25[34], c25[34]);
    FA fa610(pp[36][26], s24[34], c24[33], s25[35], c25[35]);
    FA fa611(pp[37][26], s24[35], c24[34], s25[36], c25[36]);
    FA fa612(pp[38][26], s24[36], c24[35], s25[37], c25[37]);
    FA fa613(pp[39][26], s24[37], c24[36], s25[38], c25[38]);
    FA fa614(pp[40][26], s24[38], c24[37], s25[39], c25[39]);
    FA fa615(pp[41][26], s24[39], c24[38], s25[40], c25[40]);
    FA fa616(pp[42][26], s24[40], c24[39], s25[41], c25[41]);
    FA fa617(pp[43][26], s24[41], c24[40], s25[42], c25[42]);
    FA fa618(pp[44][26], s24[42], c24[41], s25[43], c25[43]);
    FA fa619(pp[45][26], s24[43], c24[42], s25[44], c25[44]);
    FA fa620(pp[46][26], s24[44], c24[43], s25[45], c25[45]);
    FA fa621(pp[47][26], s24[45], c24[44], s25[46], c25[46]);
    FA fa622(pp[48][26], s24[46], c24[45], s25[47], c25[47]);
    FA fa623(pp[49][26], s24[47], c24[46], s25[48], c25[48]);
    FA fa624(pp[50][26], s24[48], c24[47], s25[49], c25[49]);
    FA fa625(pp[51][26], pp[52][25], c24[48], s25[50], c25[50]);

    // 26
    HA ha27(pp[26][1], pp[27][0], s26[1], c26[1]);
    FA fa626(pp[25][3], pp[26][2], s25[1], s26[2], c26[2]);
    FA fa627(pp[25][4], s25[2], c25[1], s26[3], c26[3]);
    FA fa628(pp[25][5], s25[3], c25[2], s26[4], c26[4]);
    FA fa629(pp[25][6], s25[4], c25[3], s26[5], c26[5]);
    FA fa630(pp[25][7], s25[5], c25[4], s26[6], c26[6]);
    FA fa631(pp[25][8], s25[6], c25[5], s26[7], c26[7]);
    FA fa632(pp[25][9], s25[7], c25[6], s26[8], c26[8]);
    FA fa633(pp[25][10], s25[8], c25[7], s26[9], c26[9]);
    FA fa634(pp[25][11], s25[9], c25[8], s26[10], c26[10]);
    FA fa635(pp[25][12], s25[10], c25[9], s26[11], c26[11]);
    FA fa636(pp[25][13], s25[11], c25[10], s26[12], c26[12]);
    FA fa637(pp[25][14], s25[12], c25[11], s26[13], c26[13]);
    FA fa638(pp[25][15], s25[13], c25[12], s26[14], c26[14]);
    FA fa639(pp[25][16], s25[14], c25[13], s26[15], c26[15]);
    FA fa640(pp[25][17], s25[15], c25[14], s26[16], c26[16]);
    FA fa641(pp[25][18], s25[16], c25[15], s26[17], c26[17]);
    FA fa642(pp[25][19], s25[17], c25[16], s26[18], c26[18]);
    FA fa643(pp[25][20], s25[18], c25[17], s26[19], c26[19]);
    FA fa644(pp[25][21], s25[19], c25[18], s26[20], c26[20]);
    FA fa645(pp[25][22], s25[20], c25[19], s26[21], c26[21]);
    FA fa646(pp[25][23], s25[21], c25[20], s26[22], c26[22]);
    FA fa647(pp[25][24], s25[22], c25[21], s26[23], c26[23]);
    FA fa648(pp[25][25], s25[23], c25[22], s26[24], c26[24]);
    FA fa649(pp[25][26], s25[24], c25[23], s26[25], c26[25]);
    FA fa650(pp[25][27], s25[25], c25[24], s26[26], c26[26]);
    FA fa651(pp[26][27], s25[26], c25[25], s26[27], c26[27]);
    FA fa652(pp[27][27], s25[27], c25[26], s26[28], c26[28]);
    FA fa653(pp[28][27], s25[28], c25[27], s26[29], c26[29]);
    FA fa654(pp[29][27], s25[29], c25[28], s26[30], c26[30]);
    FA fa655(pp[30][27], s25[30], c25[29], s26[31], c26[31]);
    FA fa656(pp[31][27], s25[31], c25[30], s26[32], c26[32]);
    FA fa657(pp[32][27], s25[32], c25[31], s26[33], c26[33]);
    FA fa658(pp[33][27], s25[33], c25[32], s26[34], c26[34]);
    FA fa659(pp[34][27], s25[34], c25[33], s26[35], c26[35]);
    FA fa660(pp[35][27], s25[35], c25[34], s26[36], c26[36]);
    FA fa661(pp[36][27], s25[36], c25[35], s26[37], c26[37]);
    FA fa662(pp[37][27], s25[37], c25[36], s26[38], c26[38]);
    FA fa663(pp[38][27], s25[38], c25[37], s26[39], c26[39]);
    FA fa664(pp[39][27], s25[39], c25[38], s26[40], c26[40]);
    FA fa665(pp[40][27], s25[40], c25[39], s26[41], c26[41]);
    FA fa666(pp[41][27], s25[41], c25[40], s26[42], c26[42]);
    FA fa667(pp[42][27], s25[42], c25[41], s26[43], c26[43]);
    FA fa668(pp[43][27], s25[43], c25[42], s26[44], c26[44]);
    FA fa669(pp[44][27], s25[44], c25[43], s26[45], c26[45]);
    FA fa670(pp[45][27], s25[45], c25[44], s26[46], c26[46]);
    FA fa671(pp[46][27], s25[46], c25[45], s26[47], c26[47]);
    FA fa672(pp[47][27], s25[47], c25[46], s26[48], c26[48]);
    FA fa673(pp[48][27], s25[48], c25[47], s26[49], c26[49]);
    FA fa674(pp[49][27], s25[49], c25[48], s26[50], c26[50]);
    FA fa675(pp[50][27], s25[50], c25[49], s26[51], c26[51]);
    FA fa676(pp[51][27], pp[52][26], c25[50], s26[52], c26[52]);

    // 27
    HA ha28(pp[25][1], pp[26][0], s27[1], c27[1]);
    FA fa677(pp[24][3], pp[25][2], s26[1], s27[2], c27[2]);
    FA fa678(pp[24][4], s26[2], c26[1], s27[3], c27[3]);
    FA fa679(pp[24][5], s26[3], c26[2], s27[4], c27[4]);
    FA fa680(pp[24][6], s26[4], c26[3], s27[5], c27[5]);
    FA fa681(pp[24][7], s26[5], c26[4], s27[6], c27[6]);
    FA fa682(pp[24][8], s26[6], c26[5], s27[7], c27[7]);
    FA fa683(pp[24][9], s26[7], c26[6], s27[8], c27[8]);
    FA fa684(pp[24][10], s26[8], c26[7], s27[9], c27[9]);
    FA fa685(pp[24][11], s26[9], c26[8], s27[10], c27[10]);
    FA fa686(pp[24][12], s26[10], c26[9], s27[11], c27[11]);
    FA fa687(pp[24][13], s26[11], c26[10], s27[12], c27[12]);
    FA fa688(pp[24][14], s26[12], c26[11], s27[13], c27[13]);
    FA fa689(pp[24][15], s26[13], c26[12], s27[14], c27[14]);
    FA fa690(pp[24][16], s26[14], c26[13], s27[15], c27[15]);
    FA fa691(pp[24][17], s26[15], c26[14], s27[16], c27[16]);
    FA fa692(pp[24][18], s26[16], c26[15], s27[17], c27[17]);
    FA fa693(pp[24][19], s26[17], c26[16], s27[18], c27[18]);
    FA fa694(pp[24][20], s26[18], c26[17], s27[19], c27[19]);
    FA fa695(pp[24][21], s26[19], c26[18], s27[20], c27[20]);
    FA fa696(pp[24][22], s26[20], c26[19], s27[21], c27[21]);
    FA fa697(pp[24][23], s26[21], c26[20], s27[22], c27[22]);
    FA fa698(pp[24][24], s26[22], c26[21], s27[23], c27[23]);
    FA fa699(pp[24][25], s26[23], c26[22], s27[24], c27[24]);
    FA fa700(pp[24][26], s26[24], c26[23], s27[25], c27[25]);
    FA fa701(pp[24][27], s26[25], c26[24], s27[26], c27[26]);
    FA fa702(pp[24][28], s26[26], c26[25], s27[27], c27[27]);
    FA fa703(pp[25][28], s26[27], c26[26], s27[28], c27[28]);
    FA fa704(pp[26][28], s26[28], c26[27], s27[29], c27[29]);
    FA fa705(pp[27][28], s26[29], c26[28], s27[30], c27[30]);
    FA fa706(pp[28][28], s26[30], c26[29], s27[31], c27[31]);
    FA fa707(pp[29][28], s26[31], c26[30], s27[32], c27[32]);
    FA fa708(pp[30][28], s26[32], c26[31], s27[33], c27[33]);
    FA fa709(pp[31][28], s26[33], c26[32], s27[34], c27[34]);
    FA fa710(pp[32][28], s26[34], c26[33], s27[35], c27[35]);
    FA fa711(pp[33][28], s26[35], c26[34], s27[36], c27[36]);
    FA fa712(pp[34][28], s26[36], c26[35], s27[37], c27[37]);
    FA fa713(pp[35][28], s26[37], c26[36], s27[38], c27[38]);
    FA fa714(pp[36][28], s26[38], c26[37], s27[39], c27[39]);
    FA fa715(pp[37][28], s26[39], c26[38], s27[40], c27[40]);
    FA fa716(pp[38][28], s26[40], c26[39], s27[41], c27[41]);
    FA fa717(pp[39][28], s26[41], c26[40], s27[42], c27[42]);
    FA fa718(pp[40][28], s26[42], c26[41], s27[43], c27[43]);
    FA fa719(pp[41][28], s26[43], c26[42], s27[44], c27[44]);
    FA fa720(pp[42][28], s26[44], c26[43], s27[45], c27[45]);
    FA fa721(pp[43][28], s26[45], c26[44], s27[46], c27[46]);
    FA fa722(pp[44][28], s26[46], c26[45], s27[47], c27[47]);
    FA fa723(pp[45][28], s26[47], c26[46], s27[48], c27[48]);
    FA fa724(pp[46][28], s26[48], c26[47], s27[49], c27[49]);
    FA fa725(pp[47][28], s26[49], c26[48], s27[50], c27[50]);
    FA fa726(pp[48][28], s26[50], c26[49], s27[51], c27[51]);
    FA fa727(pp[49][28], s26[51], c26[50], s27[52], c27[52]);
    FA fa728(pp[50][28], s26[52], c26[51], s27[53], c27[53]);
    FA fa729(pp[51][28], pp[52][27], c26[52], s27[54], c27[54]);

    // 28
    HA ha29(pp[24][1], pp[25][0], s28[1], c28[1]);
    FA fa730(pp[23][3], pp[24][2], s27[1], s28[2], c28[2]);
    FA fa731(pp[23][4], s27[2], c27[1], s28[3], c28[3]);
    FA fa732(pp[23][5], s27[3], c27[2], s28[4], c28[4]);
    FA fa733(pp[23][6], s27[4], c27[3], s28[5], c28[5]);
    FA fa734(pp[23][7], s27[5], c27[4], s28[6], c28[6]);
    FA fa735(pp[23][8], s27[6], c27[5], s28[7], c28[7]);
    FA fa736(pp[23][9], s27[7], c27[6], s28[8], c28[8]);
    FA fa737(pp[23][10], s27[8], c27[7], s28[9], c28[9]);
    FA fa738(pp[23][11], s27[9], c27[8], s28[10], c28[10]);
    FA fa739(pp[23][12], s27[10], c27[9], s28[11], c28[11]);
    FA fa740(pp[23][13], s27[11], c27[10], s28[12], c28[12]);
    FA fa741(pp[23][14], s27[12], c27[11], s28[13], c28[13]);
    FA fa742(pp[23][15], s27[13], c27[12], s28[14], c28[14]);
    FA fa743(pp[23][16], s27[14], c27[13], s28[15], c28[15]);
    FA fa744(pp[23][17], s27[15], c27[14], s28[16], c28[16]);
    FA fa745(pp[23][18], s27[16], c27[15], s28[17], c28[17]);
    FA fa746(pp[23][19], s27[17], c27[16], s28[18], c28[18]);
    FA fa747(pp[23][20], s27[18], c27[17], s28[19], c28[19]);
    FA fa748(pp[23][21], s27[19], c27[18], s28[20], c28[20]);
    FA fa749(pp[23][22], s27[20], c27[19], s28[21], c28[21]);
    FA fa750(pp[23][23], s27[21], c27[20], s28[22], c28[22]);
    FA fa751(pp[23][24], s27[22], c27[21], s28[23], c28[23]);
    FA fa752(pp[23][25], s27[23], c27[22], s28[24], c28[24]);
    FA fa753(pp[23][26], s27[24], c27[23], s28[25], c28[25]);
    FA fa754(pp[23][27], s27[25], c27[24], s28[26], c28[26]);
    FA fa755(pp[23][28], s27[26], c27[25], s28[27], c28[27]);
    FA fa756(pp[23][29], s27[27], c27[26], s28[28], c28[28]);
    FA fa757(pp[24][29], s27[28], c27[27], s28[29], c28[29]);
    FA fa758(pp[25][29], s27[29], c27[28], s28[30], c28[30]);
    FA fa759(pp[26][29], s27[30], c27[29], s28[31], c28[31]);
    FA fa760(pp[27][29], s27[31], c27[30], s28[32], c28[32]);
    FA fa761(pp[28][29], s27[32], c27[31], s28[33], c28[33]);
    FA fa762(pp[29][29], s27[33], c27[32], s28[34], c28[34]);
    FA fa763(pp[30][29], s27[34], c27[33], s28[35], c28[35]);
    FA fa764(pp[31][29], s27[35], c27[34], s28[36], c28[36]);
    FA fa765(pp[32][29], s27[36], c27[35], s28[37], c28[37]);
    FA fa766(pp[33][29], s27[37], c27[36], s28[38], c28[38]);
    FA fa767(pp[34][29], s27[38], c27[37], s28[39], c28[39]);
    FA fa768(pp[35][29], s27[39], c27[38], s28[40], c28[40]);
    FA fa769(pp[36][29], s27[40], c27[39], s28[41], c28[41]);
    FA fa770(pp[37][29], s27[41], c27[40], s28[42], c28[42]);
    FA fa771(pp[38][29], s27[42], c27[41], s28[43], c28[43]);
    FA fa772(pp[39][29], s27[43], c27[42], s28[44], c28[44]);
    FA fa773(pp[40][29], s27[44], c27[43], s28[45], c28[45]);
    FA fa774(pp[41][29], s27[45], c27[44], s28[46], c28[46]);
    FA fa775(pp[42][29], s27[46], c27[45], s28[47], c28[47]);
    FA fa776(pp[43][29], s27[47], c27[46], s28[48], c28[48]);
    FA fa777(pp[44][29], s27[48], c27[47], s28[49], c28[49]);
    FA fa778(pp[45][29], s27[49], c27[48], s28[50], c28[50]);
    FA fa779(pp[46][29], s27[50], c27[49], s28[51], c28[51]);
    FA fa780(pp[47][29], s27[51], c27[50], s28[52], c28[52]);
    FA fa781(pp[48][29], s27[52], c27[51], s28[53], c28[53]);
    FA fa782(pp[49][29], s27[53], c27[52], s28[54], c28[54]);
    FA fa783(pp[50][29], s27[54], c27[53], s28[55], c28[55]);
    FA fa784(pp[51][29], pp[52][28], c27[54], s28[56], c28[56]);

    // 29
    HA ha30(pp[23][1], pp[24][0], s29[1], c29[1]);
    FA fa785(pp[22][3], pp[23][2], s27[1], s29[2], c29[2]);
    FA fa786(pp[22][4], s28[2], c28[1], s29[3], c29[3]);
    FA fa787(pp[22][5], s28[3], c28[2], s29[4], c29[4]);
    FA fa788(pp[22][6], s28[4], c28[3], s29[5], c29[5]);
    FA fa789(pp[22][7], s28[5], c28[4], s29[6], c29[6]);
    FA fa790(pp[22][8], s28[6], c28[5], s29[7], c29[7]);
    FA fa791(pp[22][9], s28[7], c28[6], s29[8], c29[8]);
    FA fa792(pp[22][10], s28[8], c28[7], s29[9], c29[9]);
    FA fa793(pp[22][11], s28[9], c28[8], s29[10], c29[10]);
    FA fa794(pp[22][12], s28[10], c28[9], s29[11], c29[11]);
    FA fa795(pp[22][13], s28[11], c28[10], s29[12], c29[12]);
    FA fa796(pp[22][14], s28[12], c28[11], s29[13], c29[13]);
    FA fa797(pp[22][15], s28[13], c28[12], s29[14], c29[14]);
    FA fa798(pp[22][16], s28[14], c28[13], s29[15], c29[15]);
    FA fa799(pp[22][17], s28[15], c28[14], s29[16], c29[16]);
    FA fa800(pp[22][18], s28[16], c28[15], s29[17], c29[17]);
    FA fa801(pp[22][19], s28[17], c28[16], s29[18], c29[18]);
    FA fa802(pp[22][20], s28[18], c28[17], s29[19], c29[19]);
    FA fa803(pp[22][21], s28[19], c28[18], s29[20], c29[20]);
    FA fa804(pp[22][22], s28[20], c28[19], s29[21], c29[21]);
    FA fa805(pp[22][23], s28[21], c28[20], s29[22], c29[22]);
    FA fa806(pp[22][24], s28[22], c28[21], s29[23], c29[23]);
    FA fa807(pp[22][25], s28[23], c28[22], s29[23], c29[24]);
    FA fa808(pp[22][26], s28[24], c28[23], s29[25], c29[25]);
    FA fa809(pp[22][27], s28[25], c28[24], s29[26], c29[26]);
    FA fa810(pp[22][28], s28[26], c28[25], s29[27], c29[27]);
    FA fa811(pp[22][29], s28[27], c28[26], s29[28], c29[28]);
    FA fa812(pp[22][30], s28[28], c28[27], s29[29], c29[29]);
    FA fa813(pp[23][30], s28[29], c28[28], s29[30], c29[30]);
    FA fa814(pp[24][30], s28[30], c28[29], s29[31], c29[31]);
    FA fa815(pp[25][30], s28[31], c28[30], s29[32], c29[32]);
    FA fa816(pp[26][30], s28[32], c28[31], s29[33], c29[33]);
    FA fa817(pp[27][30], s28[33], c28[32], s29[34], c29[34]);
    FA fa818(pp[28][30], s28[34], c28[33], s29[35], c29[35]);
    FA fa819(pp[29][30], s28[35], c28[34], s29[36], c29[36]);
    FA fa820(pp[30][30], s28[36], c28[35], s29[37], c29[37]);
    FA fa821(pp[31][30], s28[37], c28[36], s29[38], c29[38]);
    FA fa822(pp[32][30], s28[38], c28[37], s29[39], c29[39]);
    FA fa823(pp[33][30], s28[39], c28[38], s29[40], c29[40]);
    FA fa824(pp[34][30], s28[40], c28[39], s29[41], c29[41]);
    FA fa825(pp[35][30], s28[41], c28[40], s29[42], c29[42]);
    FA fa826(pp[36][30], s28[42], c28[41], s29[43], c29[43]);
    FA fa827(pp[37][30], s28[43], c28[42], s29[44], c29[44]);
    FA fa828(pp[38][30], s28[44], c28[43], s29[45], c29[45]);
    FA fa829(pp[39][30], s28[45], c28[44], s29[46], c29[46]);
    FA fa830(pp[40][30], s28[46], c28[45], s29[47], c29[47]);
    FA fa831(pp[41][30], s28[47], c28[46], s29[48], c29[48]);
    FA fa832(pp[42][30], s28[48], c28[47], s29[49], c29[49]);
    FA fa833(pp[43][30], s28[49], c28[48], s29[50], c29[50]);
    FA fa834(pp[44][30], s28[50], c28[49], s29[51], c29[51]);
    FA fa835(pp[45][30], s28[51], c28[50], s29[52], c29[52]);
    FA fa836(pp[46][30], s28[52], c28[51], s29[53], c29[53]);
    FA fa837(pp[47][30], s28[53], c28[52], s29[54], c29[54]);
    FA fa838(pp[48][30], s28[54], c28[53], s29[55], c29[55]);
    FA fa839(pp[49][30], s28[55], c28[54], s29[56], c29[56]);
    FA fa840(pp[50][30], s28[56], c28[55], s29[57], c29[57]);
    FA fa841(pp[51][30], pp[52][29], c28[56], s29[58], c29[58]);

    // 30
    HA ha31(pp[22][1], pp[23][0], s30[1], c30[1]);
    FA fa842(pp[21][3], pp[22][2], s29[1], s30[2], c30[2]);
    FA fa843(pp[21][4], s29[2], c29[1], s30[3], c30[3]);
    FA fa844(pp[21][5], s29[3], c29[2], s30[4], c30[4]);
    FA fa845(pp[21][6], s29[4], c29[3], s30[5], c30[5]);
    FA fa846(pp[21][7], s29[5], c29[4], s30[6], c30[6]);
    FA fa847(pp[21][8], s29[6], c29[5], s30[7], c30[7]);
    FA fa848(pp[21][9], s29[7], c29[6], s30[8], c30[8]);
    FA fa849(pp[21][10], s29[8], c29[7], s30[9], c30[9]);
    FA fa850(pp[21][11], s29[9], c29[8], s30[10], c30[10]);
    FA fa851(pp[21][12], s29[10], c29[9], s30[11], c30[11]);
    FA fa852(pp[21][13], s29[11], c29[10], s30[12], c30[12]);
    FA fa853(pp[21][14], s29[12], c29[11], s30[13], c30[13]);
    FA fa854(pp[21][15], s29[13], c29[12], s30[14], c30[14]);
    FA fa855(pp[21][16], s29[14], c29[13], s30[15], c30[15]);
    FA fa856(pp[21][17], s29[15], c29[14], s30[16], c30[16]);
    FA fa857(pp[21][18], s29[16], c29[15], s30[17], c30[17]);
    FA fa858(pp[21][19], s29[17], c29[16], s30[18], c30[18]);
    FA fa859(pp[21][20], s29[18], c29[17], s30[19], c30[19]);
    FA fa860(pp[21][21], s29[19], c29[18], s30[20], c30[20]);
    FA fa861(pp[21][22], s29[20], c29[19], s30[21], c30[21]);
    FA fa862(pp[21][23], s29[21], c29[20], s30[22], c30[22]);
    FA fa863(pp[21][24], s29[22], c29[21], s30[23], c30[23]);
    FA fa864(pp[21][25], s29[23], c29[22], s30[24], c30[24]);
    FA fa865(pp[21][26], s29[24], c29[23], s30[25], c30[25]);
    FA fa866(pp[21][27], s29[25], c29[24], s30[26], c30[26]);
    FA fa867(pp[21][28], s29[26], c29[25], s30[27], c30[27]);
    FA fa868(pp[21][29], s29[27], c29[26], s30[28], c30[28]);
    FA fa869(pp[21][30], s29[28], c29[27], s30[29], c30[29]);
    FA fa870(pp[21][31], s29[29], c29[28], s30[30], c30[30]);
    FA fa871(pp[22][31], s29[30], c29[29], s30[31], c30[31]);
    FA fa872(pp[23][31], s29[31], c29[30], s30[32], c30[32]);
    FA fa873(pp[24][31], s29[32], c29[31], s30[33], c30[33]);
    FA fa874(pp[25][31], s29[33], c29[32], s30[34], c30[34]);
    FA fa875(pp[26][31], s29[34], c29[33], s30[35], c30[35]);
    FA fa876(pp[27][31], s29[35], c29[34], s30[36], c30[36]);
    FA fa877(pp[28][31], s29[36], c29[35], s30[37], c30[37]);
    FA fa878(pp[29][31], s29[37], c29[36], s30[38], c30[38]);
    FA fa879(pp[30][31], s29[38], c29[37], s30[39], c30[39]);
    FA fa880(pp[31][31], s29[39], c29[38], s30[40], c30[40]);
    FA fa881(pp[32][31], s29[40], c29[39], s30[41], c30[41]);
    FA fa882(pp[33][31], s29[41], c29[40], s30[42], c30[42]);
    FA fa883(pp[34][31], s29[42], c29[41], s30[43], c30[43]);
    FA fa884(pp[35][31], s29[43], c29[42], s30[44], c30[44]);
    FA fa885(pp[36][31], s29[44], c29[43], s30[45], c30[45]);
    FA fa886(pp[37][31], s29[45], c29[44], s30[46], c30[46]);
    FA fa887(pp[38][31], s29[46], c29[45], s30[47], c30[47]);
    FA fa888(pp[39][31], s29[47], c29[46], s30[48], c30[48]);
    FA fa889(pp[40][31], s29[48], c29[47], s30[49], c30[49]);
    FA fa890(pp[41][31], s29[49], c29[48], s30[50], c30[50]);
    FA fa891(pp[42][31], s29[50], c29[49], s30[51], c30[51]);
    FA fa892(pp[43][31], s29[51], c29[50], s30[52], c30[52]);
    FA fa893(pp[44][31], s29[52], c29[51], s30[53], c30[53]);
    FA fa894(pp[45][31], s29[53], c29[52], s30[54], c30[54]);
    FA fa895(pp[46][31], s29[54], c29[53], s30[55], c30[55]);
    FA fa896(pp[47][31], s29[55], c29[54], s30[56], c30[56]);
    FA fa897(pp[48][31], s29[56], c29[55], s30[57], c30[57]);
    FA fa898(pp[49][31], s29[57], c29[56], s30[58], c30[58]);
    FA fa899(pp[50][31], s29[58], c29[57], s30[59], c30[59]);
    FA fa900(pp[51][31], pp[52][30], c29[58], s30[60], c30[60]);

    // 31
    HA ha32(pp[21][1], pp[22][0], s31[1], c31[1]);
    FA fa901(pp[20][3], pp[21][2], s30[1], s31[2], c31[2]);
    FA fa902(pp[20][4], s30[2], c[30][1], s31[3], c31[3]);
    FA fa903(pp[20][5], s30[3], c[30][2], s31[4], c31[4]);
    FA fa904(pp[20][6], s30[4], c[30][3], s31[5], c31[5]);
    FA fa905(pp[20][7], s30[5], c[30][4], s31[6], c31[6]);
    FA fa906(pp[20][8], s30[6], c[30][5], s31[7], c31[7]);
    FA fa907(pp[20][9], s30[7], c[30][6], s31[8], c31[8]);
    FA fa908(pp[20][10], s30[8], c[30][7], s31[9], c31[9]);
    FA fa909(pp[20][11], s30[9], c[30][8], s31[10], c31[10]);
    FA fa910(pp[20][12], s30[10], c[30][9], s31[11], c31[11]);
    FA fa911(pp[20][13], s30[11], c[30][10], s31[12], c31[12]);
    FA fa912(pp[20][14], s30[12], c[30][11], s31[13], c31[13]);
    FA fa913(pp[20][15], s30[13], c[30][12], s31[14], c31[14]);
    FA fa914(pp[20][16], s30[14], c[30][13], s31[15], c31[15]);
    FA fa915(pp[20][17], s30[15], c[30][14], s31[16], c31[16]);
    FA fa916(pp[20][18], s30[16], c[30][15], s31[17], c31[17]);
    FA fa917(pp[20][19], s30[17], c[30][16], s31[18], c32[18]);
    FA fa918(pp[20][20], s30[18], c[30][17], s31[19], c31[19]);
    FA fa919(pp[20][21], s30[19], c[30][18], s31[20], c31[20]);
    FA fa920(pp[20][22], s30[20], c[30][19], s31[21], c31[21]);
    FA fa921(pp[20][23], s30[21], c[30][20], s31[22], c31[22]);
    FA fa922(pp[20][24], s30[22], c[30][21], s31[23], c31[23]);
    FA fa923(pp[20][25], s30[23], c[30][22], s31[24], c31[24]);
    FA fa924(pp[20][26], s30[24], c[30][23], s31[25], c31[25]);
    FA fa925(pp[20][27], s30[25], c[30][24], s31[26], c31[26]);
    FA fa926(pp[20][28], s30[26], c[30][25], s31[27], c31[27]);
    FA fa927(pp[20][29], s30[27], c[30][26], s31[28], c31[28]);
    FA fa928(pp[20][30], s30[28], c[30][27], s31[29], c31[29]);
    FA fa929(pp[20][31], s30[29], c[30][28], s31[30], c31[30]);
    FA fa930(pp[20][32], s30[30], c[30][29], s31[31], c31[31]);
    FA fa931(pp[21][32], s30[31], c[30][30], s31[32], c31[32]);
    FA fa932(pp[22][32], s30[32], c[30][31], s31[33], c31[33]);
    FA fa933(pp[23][32], s30[33], c[30][32], s31[34], c31[34]);
    FA fa934(pp[24][32], s30[34], c[30][33], s31[35], c31[35]);
    FA fa935(pp[25][32], s30[35], c[30][34], s31[36], c31[36]);
    FA fa936(pp[26][32], s30[36], c[30][35], s31[37], c31[37]);
    FA fa937(pp[27][32], s30[37], c[30][36], s31[38], c31[38]);
    FA fa938(pp[28][32], s30[38], c[30][37], s31[39], c31[39]);
    FA fa939(pp[29][32], s30[39], c[30][38], s31[40], c31[40]);
    FA fa940(pp[30][32], s30[40], c[30][39], s31[41], c31[41]);
    FA fa941(pp[31][32], s30[41], c[30][40], s31[42], c31[42]);
    FA fa942(pp[32][32], s30[42], c[30][41], s31[43], c31[43]);
    FA fa943(pp[33][32], s30[43], c[30][42], s31[44], c31[44]);
    FA fa944(pp[34][32], s30[44], c[30][43], s31[45], c31[45]);
    FA fa945(pp[35][32], s30[45], c[30][44], s31[46], c31[46]);
    FA fa946(pp[36][32], s30[46], c[30][45], s31[47], c31[47]);
    FA fa947(pp[37][32], s30[47], c[30][46], s31[48], c31[48]);
    FA fa948(pp[38][32], s30[48], c[30][47], s31[49], c31[49]);
    FA fa949(pp[39][32], s30[49], c[30][48], s31[50], c31[50]);
    FA fa950(pp[40][32], s30[50], c[30][49], s31[51], c31[51]);
    FA fa951(pp[41][32], s30[51], c[30][50], s31[52], c31[52]);
    FA fa952(pp[42][32], s30[52], c[30][51], s31[53], c31[53]);
    FA fa953(pp[43][32], s30[53], c[30][52], s31[54], c31[54]);
    FA fa954(pp[44][32], s30[54], c[30][53], s31[55], c31[55]);
    FA fa955(pp[45][32], s30[55], c[30][54], s31[56], c31[56]);
    FA fa956(pp[46][32], s30[56], c[30][55], s31[57], c31[57]);
    FA fa957(pp[47][32], s30[57], c[30][56], s31[58], c31[58]);
    FA fa958(pp[48][32], s30[58], c[30][57], s31[59], c31[59]);
    FA fa959(pp[49][32], s30[59], c[30][58], s31[60], c31[60]);
    FA fa960(pp[50][32], s30[60], c[30][59], s31[61], c31[61]);
    FA fa961(pp[51][32], pp[52][31], c[30][60], s31[62], c31[62]);

    // 32
    HA ha33(pp[20][1], pp[21][0], s32[1], c32[1]);
    FA fa962(pp[19][3], pp[20][2], s31[1], s32[2], c32[2]);
    FA fa963(pp[19][4], s31[2], c31[1], s32[3], c32[3]);
    FA fa964(pp[19][5], s31[3], c31[2], s32[4], c32[4]);
    FA fa965(pp[19][6], s31[4], c31[3], s32[5], c32[5]);
    FA fa966(pp[19][7], s31[5], c31[4], s32[6], c32[6]);
    FA fa967(pp[19][8], s31[6], c31[5], s32[7], c32[7]);
    FA fa968(pp[19][9], s31[7], c31[6], s32[8], c32[8]);
    FA fa969(pp[19][10], s31[8], c31[7], s32[9], c32[9]);
    FA fa970(pp[19][11], s31[9], c31[8], s32[10], c32[10]);
    FA fa971(pp[19][12], s31[10], c31[9], s32[11], c32[11]);
    FA fa972(pp[19][13], s31[11], c31[10], s32[12], c32[12]);
    FA fa973(pp[19][14], s31[12], c31[11], s32[13], c32[13]);
    FA fa974(pp[19][15], s31[13], c31[12], s32[14], c32[14]);
    FA fa975(pp[19][16], s31[14], c31[13], s32[15], c32[15]);
    FA fa976(pp[19][17], s31[15], c31[14], s32[16], c32[16]);
    FA fa977(pp[19][18], s31[16], c31[15], s32[17], c32[17]);
    FA fa978(pp[19][19], s31[17], c31[16], s32[18], c32[18]);
    FA fa979(pp[19][20], s31[18], c31[17], s32[19], c32[19]);
    FA fa980(pp[19][21], s31[19], c31[18], s32[20], c32[20]);
    FA fa981(pp[19][22], s31[20], c31[19], s32[21], c32[21]);
    FA fa982(pp[19][23], s31[21], c31[20], s32[22], c32[22]);
    FA fa983(pp[19][24], s31[22], c31[21], s32[23], c32[23]);
    FA fa984(pp[19][25], s31[23], c31[22], s32[24], c32[24]);
    FA fa985(pp[19][26], s31[24], c31[23], s32[25], c32[25]);
    FA fa986(pp[19][27], s31[25], c31[24], s32[26], c32[26]);
    FA fa987(pp[19][28], s31[26], c31[25], s32[27], c32[27]);
    FA fa988(pp[19][29], s31[27], c31[26], s32[28], c32[28]);
    FA fa989(pp[19][30], s31[28], c31[27], s32[29], c32[29]);
    FA fa990(pp[19][31], s31[29], c31[28], s32[30], c32[30]);
    FA fa991(pp[19][32], s31[30], c31[29], s32[31], c32[31]);
    FA fa992(pp[19][33], s31[31], c31[30], s32[32], c32[32]);
    FA fa993(pp[20][33], s31[32], c31[31], s32[33], c32[33]);
    FA fa994(pp[21][33], s31[33], c31[32], s32[34], c32[34]);
    FA fa995(pp[22][33], s31[34], c31[33], s32[35], c32[35]);
    FA fa996(pp[23][33], s31[35], c31[34], s32[36], c32[36]);
    FA fa997(pp[24][33], s31[36], c31[35], s32[37], c32[37]);
    FA fa998(pp[25][33], s31[37], c31[36], s32[38], c32[38]);
    FA fa999(pp[26][33], s31[38], c31[37], s32[39], c32[39]);
    FA fa1000(pp[27][33], s31[39], c31[38], s32[40], c32[40]);
    FA fa1001(pp[28][33], s31[40], c31[39], s32[41], c32[41]);
    FA fa1002(pp[29][33], s31[41], c31[40], s32[42], c32[42]);
    FA fa1003(pp[30][33], s31[42], c31[41], s32[43], c32[43]);
    FA fa1004(pp[31][33], s31[43], c31[42], s32[44], c32[44]);
    FA fa1005(pp[32][33], s31[44], c31[43], s32[45], c32[45]);
    FA fa1006(pp[33][33], s31[45], c31[44], s32[46], c32[46]);
    FA fa1007(pp[34][33], s31[46], c31[45], s32[47], c32[47]);
    FA fa1008(pp[35][33], s31[47], c31[46], s32[48], c32[48]);
    FA fa1009(pp[36][33], s31[48], c31[47], s32[49], c32[49]);
    FA fa1010(pp[37][33], s31[49], c31[48], s32[50], c32[50]);
    FA fa1011(pp[38][33], s31[50], c31[49], s32[51], c32[51]);
    FA fa1012(pp[39][33], s31[51], c31[50], s32[52], c32[52]);
    FA fa1013(pp[40][33], s31[52], c31[51], s32[53], c32[53]);
    FA fa1014(pp[41][33], s31[53], c31[52], s32[54], c32[54]);
    FA fa1015(pp[42][33], s31[54], c31[53], s32[55], c32[55]);
    FA fa1016(pp[43][33], s31[55], c31[54], s32[56], c32[56]);
    FA fa1017(pp[44][33], s31[56], c31[55], s32[57], c32[57]);
    FA fa1018(pp[45][33], s31[57], c31[56], s32[58], c32[58]);
    FA fa1019(pp[46][33], s31[58], c31[57], s32[59], c32[59]);
    FA fa1020(pp[47][33], s31[59], c31[58], s32[60], c32[60]);
    FA fa1021(pp[48][33], s31[60], c31[59], s32[61], c32[61]);
    FA fa1022(pp[49][33], s31[61], c31[60], s32[62], c32[62]);
    FA fa1023(pp[50][33], s31[62], c31[61], s32[63], c32[63]);
    FA fa1024(pp[51][33], pp[52][32], c31[62], s32[64], c32[64]);

    // 33
    HA ha31(pp[19][1], pp[20][0], s33[1], c33[1]);
    FA fa1025(pp[18][3], pp[19][2], s32[1], s33[2], c33[2]);
    FA fa1026();
    FA fa1027();
    FA fa1028();
    FA fa1029();
    FA fa1030();
    FA fa1031();
    FA fa1032();
    FA fa1033();
    FA fa1034();
    FA fa1035();
    FA fa1036();
    FA fa1037();
    FA fa1038();
    FA fa1039();
    FA fa1040();
    FA fa1041();
    FA fa1042();
    FA fa1043();
    FA fa1044();
    FA fa1045();
    FA fa1046();
    FA fa1047();
    FA fa1048();
    FA fa1049();
    FA fa1050();
    FA fa1051();
    FA fa1052();
    FA fa1053();
    FA fa1054();
    FA fa1055();
    FA fa1056();
    FA fa1057();
    FA fa1058();
    FA fa1059();
    FA fa1060();
    FA fa1061();
    FA fa1062();
    FA fa1063();
    FA fa1064();
    FA fa1065();
    FA fa1066();
    FA fa1067();
    FA fa1068();
    FA fa1069();
    FA fa1070();
    FA fa1071();
    FA fa1072();
    FA fa1073();
    FA fa1074();
    FA fa1075();
    FA fa1076();
    FA fa1077();
    FA fa1078();
    FA fa1079();
    FA fa1080();
    FA fa1081();
    FA fa1082();
    FA fa1083();
    FA fa1084();
    FA fa1085();
    FA fa1086();
    FA fa1087();
    FA fa1088();
    FA fa1089();
    FA fa1090();
    FA fa1091();
    FA fa1092();
    FA fa1093();
    FA fa1094();
    FA fa1095();
    FA fa1096();
    FA fa1097();
    FA fa1098();
    FA fa1099();
    FA fa1100();
    FA fa1101();
    FA fa1102();
    FA fa1103();
    FA fa1104();
    FA fa1105();
    FA fa1106();
    FA fa1107();
    FA fa1108();
    FA fa1109();
    FA fa1110();
    FA fa1111();
    FA fa1112();
    FA fa1113();
    FA fa1114();
    FA fa1115();
    FA fa1116();
    FA fa1117();
    FA fa1118();
    FA fa1119();
    FA fa1120();
    FA fa1121();
    FA fa1122();
    FA fa1123();
    FA fa1124();
    FA fa1125();
    FA fa1126();
    FA fa1127();
    FA fa1128();
    FA fa1129();
    FA fa1130();
    FA fa1131();
    FA fa1132();
    FA fa1133();
    FA fa1134();
    FA fa1135();
    FA fa1136();
    FA fa1137();
    FA fa1138();
    FA fa1139();
    FA fa1140();
    FA fa1141();
    FA fa1142();
    FA fa1143();
    FA fa1144();
    FA fa1145();
    FA fa1146();
    FA fa1147();
    FA fa1148();
    FA fa1149();
    FA fa1150();
    FA fa1151();
    FA fa1152();
    FA fa1153();
    FA fa1154();
    FA fa1155();
    FA fa1156();
    FA fa1157();
    FA fa1158();
    FA fa1159();
    FA fa1160();
    FA fa1161();
    FA fa1162();
    FA fa1163();
    FA fa1164();
    FA fa1165();
    FA fa1166();
    FA fa1167();
    FA fa1168();
    FA fa1169();
    FA fa1170();
    FA fa1171();
    FA fa1172();
    FA fa1173();
    FA fa1174();
    FA fa1175();
    FA fa1176();
    FA fa1177();
    FA fa1178();
    FA fa1179();
    FA fa1180();
    FA fa1181();
    FA fa1182();
    FA fa1183();
    FA fa1184();
    FA fa1185();
    FA fa1186();
    FA fa1187();
    FA fa1188();
    FA fa1189();
    FA fa1190();
    FA fa1191();
    FA fa1192();
    FA fa1193();
    FA fa1194();
    FA fa1195();
    FA fa1196();
    FA fa1197();
    FA fa1198();
    FA fa1199();
    FA fa1200();
    FA fa1201();
    FA fa1202();
    FA fa1203();
    FA fa1204();
    FA fa1205();
    FA fa1206();
    FA fa1207();
    FA fa1208();
    FA fa1209();
    FA fa1210();
    FA fa1211();
    FA fa1212();
    FA fa1213();
    FA fa1214();
    FA fa1215();
    FA fa1216();
    FA fa1217();
    FA fa1218();
    FA fa1219();
    FA fa1220();
    FA fa1221();
    FA fa1222();
    FA fa1223();
    FA fa1224();
    FA fa1225();
    FA fa1226();
    FA fa1227();
    FA fa1228();
    FA fa1229();
    FA fa1230();
    FA fa1231();
    FA fa1232();
    FA fa1233();
    FA fa1234();
    FA fa1235();
    FA fa1236();
    FA fa1237();
    FA fa1238();
    FA fa1239();
    FA fa1240();
    FA fa1241();
    FA fa1242();
    FA fa1243();
    FA fa1244();
    FA fa1245();
    FA fa1246();
    FA fa1247();
    FA fa1248();
    FA fa1249();
    FA fa1250();
    FA fa1251();
    FA fa1252();
    FA fa1253();
    FA fa1254();
    FA fa1255();
    FA fa1256();
    FA fa1257();
    FA fa1258();
    FA fa1259();
    FA fa1260();
    FA fa1261();
    FA fa1262();
    FA fa1263();
    FA fa1264();
    FA fa1265();
    FA fa1266();
    FA fa1267();
    FA fa1268();
    FA fa1269();
    FA fa1270();
    FA fa1271();
    FA fa1272();
    FA fa1273();
    FA fa1274();
    FA fa1275();
    FA fa1276();
    FA fa1277();
    FA fa1278();
    FA fa1279();
    FA fa1280();
    FA fa1281();
    FA fa1282();
    FA fa1283();
    FA fa1284();
    FA fa1285();
    FA fa1286();
    FA fa1287();
    FA fa1288();
    FA fa1289();
    FA fa1290();
    FA fa1291();
    FA fa1292();
    FA fa1293();
    FA fa1294();
    FA fa1295();
    FA fa1296();
    FA fa1297();
    FA fa1298();
    FA fa1299();
    FA fa1300();
    FA fa1301();
    FA fa1302();
    FA fa1303();
    FA fa1304();
    FA fa1305();
    FA fa1306();
    FA fa1307();
    FA fa1308();
    FA fa1309();
    FA fa1310();
    FA fa1311();
    FA fa1312();
    FA fa1313();
    FA fa1314();
    FA fa1315();
    FA fa1316();
    FA fa1317();
    FA fa1318();
    FA fa1319();
    FA fa1320();
    FA fa1321();
    FA fa1322();
    FA fa1323();
    FA fa1324();
    FA fa1325();
    FA fa1326();
    FA fa1327();
    FA fa1328();
    FA fa1329();
    FA fa1330();
    FA fa1331();
    FA fa1332();
    FA fa1333();
    FA fa1334();
    FA fa1335();
    FA fa1336();
    FA fa1337();
    FA fa1338();
    FA fa1339();
    FA fa1340();
    FA fa1341();
    FA fa1342();
    FA fa1343();
    FA fa1344();
    FA fa1345();
    FA fa1346();
    FA fa1347();
    FA fa1348();
    FA fa1349();
    FA fa1350();
    FA fa1351();
    FA fa1352();
    FA fa1353();
    FA fa1354();
    FA fa1355();
    FA fa1356();
    FA fa1357();
    FA fa1358();
    FA fa1359();
    FA fa1360();
    FA fa1361();
    FA fa1362();
    FA fa1363();
    FA fa1364();
    FA fa1365();
    FA fa1366();
    FA fa1367();
    FA fa1368();
    FA fa1369();
    FA fa1370();
    FA fa1371();
    FA fa1372();
    FA fa1373();
    FA fa1374();
    FA fa1375();
    FA fa1376();
    FA fa1377();
    FA fa1378();
    FA fa1379();
    FA fa1380();
    FA fa1381();
    FA fa1382();
    FA fa1383();
    FA fa1384();
    FA fa1385();
    FA fa1386();
    FA fa1387();
    FA fa1388();
    FA fa1389();
    FA fa1390();
    FA fa1391();
    FA fa1392();
    FA fa1393();
    FA fa1394();
    FA fa1395();
    FA fa1396();
    FA fa1397();
    FA fa1398();
    FA fa1399();
    FA fa1400();
    FA fa1401();
    FA fa1402();
    FA fa1403();
    FA fa1404();
    FA fa1405();
    FA fa1406();
    FA fa1407();
    FA fa1408();
    FA fa1409();
    FA fa1410();
    FA fa1411();
    FA fa1412();
    FA fa1413();
    FA fa1414();
    FA fa1415();
    FA fa1416();
    FA fa1417();
    FA fa1418();
    FA fa1419();
    FA fa1420();
    FA fa1421();
    FA fa1422();
    FA fa1423();
    FA fa1424();
    FA fa1425();
    FA fa1426();
    FA fa1427();
    FA fa1428();
    FA fa1429();
    FA fa1430();
    FA fa1431();
    FA fa1432();
    FA fa1433();
    FA fa1434();
    FA fa1435();
    FA fa1436();
    FA fa1437();
    FA fa1438();
    FA fa1439();
    FA fa1440();
    FA fa1441();
    FA fa1442();
    FA fa1443();
    FA fa1444();
    FA fa1445();
    FA fa1446();
    FA fa1447();
    FA fa1448();
    FA fa1449();
    FA fa1450();
    FA fa1451();
    FA fa1452();
    FA fa1453();
    FA fa1454();
    FA fa1455();
    FA fa1456();
    FA fa1457();
    FA fa1458();
    FA fa1459();
    FA fa1460();
    FA fa1461();
    FA fa1462();
    FA fa1463();
    FA fa1464();
    FA fa1465();
    FA fa1466();
    FA fa1467();
    FA fa1468();
    FA fa1469();
    FA fa1470();
    FA fa1471();
    FA fa1472();
    FA fa1473();
    FA fa1474();
    FA fa1475();
    FA fa1476();
    FA fa1477();
    FA fa1478();
    FA fa1479();
    FA fa1480();
    FA fa1481();
    FA fa1482();
    FA fa1483();
    FA fa1484();
    FA fa1485();
    FA fa1486();
    FA fa1487();
    FA fa1488();
    FA fa1489();
    FA fa1490();
    FA fa1491();
    FA fa1492();
    FA fa1493();
    FA fa1494();
    FA fa1495();
    FA fa1496();
    FA fa1497();
    FA fa1498();
    FA fa1499();
    FA fa1500();
    FA fa1501();
    FA fa1502();
    FA fa1503();
    FA fa1504();
    FA fa1505();
    FA fa1506();
    FA fa1507();
    FA fa1508();
    FA fa1509();
    FA fa1510();
    FA fa1511();
    FA fa1512();
    FA fa1513();
    FA fa1514();
    FA fa1515();
    FA fa1516();
    FA fa1517();
    FA fa1518();
    FA fa1519();
    FA fa1520();
    FA fa1521();
    FA fa1522();
    FA fa1523();
    FA fa1524();
    FA fa1525();
    FA fa1526();
    FA fa1527();
    FA fa1528();
    FA fa1529();
    FA fa1530();
    FA fa1531();
    FA fa1532();
    FA fa1533();
    FA fa1534();
    FA fa1535();
    FA fa1536();
    FA fa1537();
    FA fa1538();
    FA fa1539();
    FA fa1540();
    FA fa1541();
    FA fa1542();
    FA fa1543();
    FA fa1544();
    FA fa1545();
    FA fa1546();
    FA fa1547();
    FA fa1548();
    FA fa1549();
    FA fa1550();
    FA fa1551();
    FA fa1552();
    FA fa1553();
    FA fa1554();
    FA fa1555();
    FA fa1556();
    FA fa1557();
    FA fa1558();
    FA fa1559();
    FA fa1560();
    FA fa1561();
    FA fa1562();
    FA fa1563();
    FA fa1564();
    FA fa1565();
    FA fa1566();
    FA fa1567();
    FA fa1568();
    FA fa1569();
    FA fa1570();
    FA fa1571();
    FA fa1572();
    FA fa1573();
    FA fa1574();
    FA fa1575();
    FA fa1576();
    FA fa1577();
    FA fa1578();
    FA fa1579();
    FA fa1580();
    FA fa1581();
    FA fa1582();
    FA fa1583();
    FA fa1584();
    FA fa1585();
    FA fa1586();
    FA fa1587();
    FA fa1588();
    FA fa1589();
    FA fa1590();
    FA fa1591();
    FA fa1592();
    FA fa1593();
    FA fa1594();
    FA fa1595();
    FA fa1596();
    FA fa1597();
    FA fa1598();
    FA fa1599();
    FA fa1600();



    


    assign pro = pp[52]; //pp[51] gives ma&53{mb[51]}; pp[51][51] gives 51st bit in pp[51]
endmodule


// 0000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000
// 0000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000
// 0000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000


// Main module 
module FP_MUL(a, b, out, out1, out2, out3, out4, out5, out6, out7);
// module FP_MUL (a, b, out);
    input[63:0] a, b; 
    // output[63:0] out;
  
    output[52:0] out, out1;
    output[52:0] out4;
    output out2, out3, out5;
    output[10:0] out6;
    output[51:0] out7;

    wire[63:0] new_a, new_b;        // Variable for new inputs that r used after swapping small one to b 
    wire sa, sb;                    // Variables for storing signs of original inputs 
    wire[10:0] ea, eb;              // Variables for storing expo of original inputs 
    wire[52:0] ma, mb;              // Variables for storing mantissa of original inputs

    wire[52:0] pro;

    // Declaring output indvivdual variables 
    wire sr_ini;
    reg sr; 
    reg[10:0] er; 
    reg[51:0] mr; 
    reg[1:0] temp;

    wire[10:0] zeroes, ones;
    wire[52:0] zeroes1, ones1;

    assign zeroes = 11'b00000000000;
    assign zeroes1 = 52'b0000000000000000000000000000000000000000000000000000;
    assign ones = 11'b11111111111;
    assign ones1 = 52'b1111111111111111111111111111111111111111111111111111;

    // Assigning the components to inputs to individual variables. Added one before mantissa that is 1 before decimal 
    assign sa = a[63]; 
    assign ea = a[62: 52]; 
    assign ma = {1'b1,a[51:0]};
    assign sb = b[63]; 
    assign eb = b[62: 52]; 
    assign mb = {1'b1,b[51:0]};

    always @(a, b) begin
        if ((ea[10:0]==ones & ma[51:0]==zeroes1) | (eb[10:0]==ones & mb[51:0]==zeroes1)) begin
            // Either number is zero
            temp = 2'b00;
        end
        else if ((ea[10:0]==zeroes & ma[51:0]==zeroes1) | (eb[10:0]==zeroes & mb[51:0]==zeroes1)) begin
            // Either number is INF
            temp = 2'b01;
        end
        else begin
            temp = 2'b10;
        end
    end

    MUL_MANT mul_mant1(ma, mb, pro);


    always @(*) begin
        if (temp==2'b00) begin
            sr = 0;
            er = ones;
            mr = 0;
        end
        else if(temp==2'b01)begin
            sr = 0;
            er = zeroes;
            mr = 0;
        end
    end


    assign out  = ma;
    assign out1 = mb;
    assign out2 = sa;
    assign out3 = sb;
    assign out4 = pro;
    assign out5 = sr;
    assign out6 = er;
    // assign out6 = er;
    assign out7 = mr;
    // assign out7 = 0;
endmodule






module FP_MUL_TB;
    reg[63:0] a, b;

    wire[52:0] res, res1;
    wire[52:0] res4;
    wire res2, res3, res5;
    wire[10:0] res6;
    wire[51:0] res7;

    // wire[63:0] out;

    FP_MUL fp_mul1(a, b, res, res1, res2, res3, res4, res5, res6, res7);
    // FP_MUL fp_mul1(a, b, out);

    initial begin
        // a=1.5; b=1.0000000000000002
        #0 a=64'b0011111111111000000000000000000000000000000000000000000000000000; b=64'b0011111111110000000000000000000000000000000000000000000000000001;
        
        // a=1.5; b=-3
        #10 a=64'b0011111111111000000000000000000000000000000000000000000000000000; b=64'b1100000000001000000000000000000000000000000000000000000000000000;

        // a=1; b=-2
        #10 a=64'b0011111111110000000000000000000000000000000000000000000000000000; b=64'b1100000000000000000000000000000000000000000000000000000000000000;

        // a=0
        #10 a=64'b0000000000000000000000000000000000000000000000000000000000000000; b=64'b1100000000001000000000000000000000000000000000000000000000000000;

        // b=-0
        #10 a=64'b0011111111111000000000000000000000000000000000000000000000000000; b=64'b1000000000000000000000000000000000000000000000000000000000000000;

        // a=INF
        #10 a=64'b0111111111110000000000000000000000000000000000000000000000000000; b=64'b1100000000001000000000000000000000000000000000000000000000000000;

        // b=-INF
        #10 a=64'b0011111111111000000000000000000000000000000000000000000000000000; b=64'b1111111111110000000000000000000000000000000000000000000000000000;
    end

    initial begin
        // $monitor(" a=%b b=%b Pro=%b", a, b, out);
        $monitor("%d: a=%b b=%b ma=%b mb=%b sa=%b sb=%b sum=%b sign=%b exp=%b man=%b", $time, a, b, res, res1, res2, res3, res4, res5, res6, res7);
    end


endmodule