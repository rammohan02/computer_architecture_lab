


module LOGIC_UNIT_TB ;
    reg[63:0] in1, in2;

    reg[2:0] sel;

    wire[63:0] out;

    LOGIC_UNIT logic_unit1(in1, in2, sel, out);

    initial begin
        #0 in1=64'b0010010101010110110110111010000100010001100100010100010001011010;in2=64'b0111000110000110100110000110000111011110110111100111001110111011; sel=3'b000;

        // #10 in1=64'b1101100111101111000101001000101001011011101100001110001100001100;                                                       in2=64'b0111010010010101010000111011110010111001110001100000000001001000; sel=3'b001;

        
        // #10 in1=64'b1111111111111111111111111111111111111111111111111111111111111111;                                                       in2=64'b1111111111111111111111111111111111111111111111111111111111111111; sel=3'b010;
        
        #10 sel=3'b001;
        #10 sel=3'b010;
        #10 sel=3'b011;
        #10 sel=3'b100;
        #10 sel=3'b101;
        #10 sel=3'b110;
        #10 sel=3'b111;

        #10;
    end

    initial begin
        $monitor("in1=%b \nin2=%b \nsel=%b \nout=%b\n", in1, in2, sel, out);
        $dumpfile("logic_unit.vcd");
        $dumpvars(0, logic_unit1);
    end


endmodule