
// Test bench
module WALLACE_TB;
    reg[63:0] a, b;

    wire[127:0] out;
    wire carry;

    WALLACE wallace1(a, b, out, carry);

    initial begin
        #0 a=64'b0000000000000000000000000000000000000000000000000000000000001000;                                                      b=64'b0000000000000000000000000000000000000000000000000000000000000100;

        #10 a=64'b0000000000000000000000000000000000000000000000000000000000001111;                                                      b=64'b0000000000000000000000000000000000000000000000000000000000001111;

        #10 a=64'b0011110100111001000101101110101010110001000000001011000011110010; b=64'b1001010011111101010011000101001100111101111000100111011111111001; 
    end

    initial begin
        $monitor("\n in1=%b, in2=%b, pro=%b", a, b, out);
        $dumpfile("wallace.vcd");
        $dumpvars(0, wallace1);
    end
endmodule